VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO trng_wb_wrapper
  CLASS BLOCK ;
  FOREIGN trng_wb_wrapper ;
  ORIGIN 0.000 0.000 ;
  SIZE 200.000 BY 300.000 ;
  PIN rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 146.240 200.000 146.840 ;
    END
  END rst_i
  PIN trng_buffer_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.950 296.000 42.230 300.000 ;
    END
  END trng_buffer_o[0]
  PIN trng_buffer_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 81.640 4.000 82.240 ;
    END
  END trng_buffer_o[10]
  PIN trng_buffer_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.130 296.000 103.410 300.000 ;
    END
  END trng_buffer_o[11]
  PIN trng_buffer_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 210.840 4.000 211.440 ;
    END
  END trng_buffer_o[12]
  PIN trng_buffer_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.240 4.000 27.840 ;
    END
  END trng_buffer_o[13]
  PIN trng_buffer_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 163.240 4.000 163.840 ;
    END
  END trng_buffer_o[14]
  PIN trng_buffer_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 108.840 4.000 109.440 ;
    END
  END trng_buffer_o[15]
  PIN trng_buffer_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.290 296.000 32.570 300.000 ;
    END
  END trng_buffer_o[16]
  PIN trng_buffer_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.050 0.000 58.330 4.000 ;
    END
  END trng_buffer_o[17]
  PIN trng_buffer_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.990 0.000 145.270 4.000 ;
    END
  END trng_buffer_o[18]
  PIN trng_buffer_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.750 296.000 171.030 300.000 ;
    END
  END trng_buffer_o[19]
  PIN trng_buffer_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 34.040 200.000 34.640 ;
    END
  END trng_buffer_o[1]
  PIN trng_buffer_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 272.040 200.000 272.640 ;
    END
  END trng_buffer_o[20]
  PIN trng_buffer_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.750 0.000 171.030 4.000 ;
    END
  END trng_buffer_o[21]
  PIN trng_buffer_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 61.240 200.000 61.840 ;
    END
  END trng_buffer_o[22]
  PIN trng_buffer_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 255.040 200.000 255.640 ;
    END
  END trng_buffer_o[23]
  PIN trng_buffer_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.370 296.000 77.650 300.000 ;
    END
  END trng_buffer_o[24]
  PIN trng_buffer_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 292.440 4.000 293.040 ;
    END
  END trng_buffer_o[25]
  PIN trng_buffer_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 282.240 200.000 282.840 ;
    END
  END trng_buffer_o[26]
  PIN trng_buffer_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.190 296.000 16.470 300.000 ;
    END
  END trng_buffer_o[27]
  PIN trng_buffer_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 153.040 4.000 153.640 ;
    END
  END trng_buffer_o[28]
  PIN trng_buffer_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 27.240 200.000 27.840 ;
    END
  END trng_buffer_o[29]
  PIN trng_buffer_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.610 0.000 51.890 4.000 ;
    END
  END trng_buffer_o[2]
  PIN trng_buffer_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.810 296.000 84.090 300.000 ;
    END
  END trng_buffer_o[30]
  PIN trng_buffer_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 0.040 200.000 0.640 ;
    END
  END trng_buffer_o[31]
  PIN trng_buffer_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.290 0.000 32.570 4.000 ;
    END
  END trng_buffer_o[3]
  PIN trng_buffer_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.050 296.000 58.330 300.000 ;
    END
  END trng_buffer_o[4]
  PIN trng_buffer_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 108.840 200.000 109.440 ;
    END
  END trng_buffer_o[5]
  PIN trng_buffer_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 6.840 4.000 7.440 ;
    END
  END trng_buffer_o[6]
  PIN trng_buffer_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 244.840 4.000 245.440 ;
    END
  END trng_buffer_o[7]
  PIN trng_buffer_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 180.240 4.000 180.840 ;
    END
  END trng_buffer_o[8]
  PIN trng_buffer_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 154.650 296.000 154.930 300.000 ;
    END
  END trng_buffer_o[9]
  PIN trng_valid_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.230 0.000 119.510 4.000 ;
    END
  END trng_valid_o
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 288.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 288.560 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 288.560 ;
    END
  END vssd1
  PIN wb_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 119.040 200.000 119.640 ;
    END
  END wb_ack_o
  PIN wb_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 265.240 200.000 265.840 ;
    END
  END wb_adr_i[0]
  PIN wb_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 238.040 200.000 238.640 ;
    END
  END wb_adr_i[1]
  PIN wb_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 217.640 200.000 218.240 ;
    END
  END wb_adr_i[2]
  PIN wb_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 210.840 200.000 211.440 ;
    END
  END wb_adr_i[3]
  PIN wb_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.130 0.000 103.410 4.000 ;
    END
  END wb_adr_i[4]
  PIN wb_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.040 4.000 17.640 ;
    END
  END wb_adr_i[5]
  PIN wb_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 292.440 200.000 293.040 ;
    END
  END wb_adr_i[6]
  PIN wb_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 173.440 4.000 174.040 ;
    END
  END wb_adr_i[7]
  PIN wb_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.710 296.000 67.990 300.000 ;
    END
  END wb_adr_i[8]
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 173.440 200.000 174.040 ;
    END
  END wb_clk_i
  PIN wb_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 180.240 200.000 180.840 ;
    END
  END wb_cyc_i
  PIN wb_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.850 296.000 26.130 300.000 ;
    END
  END wb_dat_i[0]
  PIN wb_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.470 296.000 93.750 300.000 ;
    END
  END wb_dat_i[10]
  PIN wb_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.410 296.000 180.690 300.000 ;
    END
  END wb_dat_i[11]
  PIN wb_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.710 0.000 67.990 4.000 ;
    END
  END wb_dat_i[12]
  PIN wb_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 98.640 200.000 99.240 ;
    END
  END wb_dat_i[13]
  PIN wb_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 71.440 200.000 72.040 ;
    END
  END wb_dat_i[14]
  PIN wb_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 125.840 4.000 126.440 ;
    END
  END wb_dat_i[15]
  PIN wb_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.190 0.000 16.470 4.000 ;
    END
  END wb_dat_i[16]
  PIN wb_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 17.040 200.000 17.640 ;
    END
  END wb_dat_i[17]
  PIN wb_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 88.440 200.000 89.040 ;
    END
  END wb_dat_i[18]
  PIN wb_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.510 296.000 196.790 300.000 ;
    END
  END wb_dat_i[19]
  PIN wb_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 61.240 4.000 61.840 ;
    END
  END wb_dat_i[1]
  PIN wb_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.070 0.000 190.350 4.000 ;
    END
  END wb_dat_i[20]
  PIN wb_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.470 0.000 93.750 4.000 ;
    END
  END wb_dat_i[21]
  PIN wb_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 125.840 200.000 126.440 ;
    END
  END wb_dat_i[22]
  PIN wb_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.530 296.000 6.810 300.000 ;
    END
  END wb_dat_i[23]
  PIN wb_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 200.640 4.000 201.240 ;
    END
  END wb_dat_i[24]
  PIN wb_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 54.440 200.000 55.040 ;
    END
  END wb_dat_i[25]
  PIN wb_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 238.040 4.000 238.640 ;
    END
  END wb_dat_i[26]
  PIN wb_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.240 4.000 44.840 ;
    END
  END wb_dat_i[27]
  PIN wb_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.230 296.000 119.510 300.000 ;
    END
  END wb_dat_i[28]
  PIN wb_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.040 4.000 34.640 ;
    END
  END wb_dat_i[29]
  PIN wb_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.850 0.000 26.130 4.000 ;
    END
  END wb_dat_i[2]
  PIN wb_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.370 0.000 77.650 4.000 ;
    END
  END wb_dat_i[30]
  PIN wb_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 44.240 200.000 44.840 ;
    END
  END wb_dat_i[31]
  PIN wb_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 190.440 200.000 191.040 ;
    END
  END wb_dat_i[3]
  PIN wb_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 136.040 200.000 136.640 ;
    END
  END wb_dat_i[4]
  PIN wb_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.410 0.000 180.690 4.000 ;
    END
  END wb_dat_i[5]
  PIN wb_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 190.440 4.000 191.040 ;
    END
  END wb_dat_i[6]
  PIN wb_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 146.240 4.000 146.840 ;
    END
  END wb_dat_i[7]
  PIN wb_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 136.040 4.000 136.640 ;
    END
  END wb_dat_i[8]
  PIN wb_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 153.040 200.000 153.640 ;
    END
  END wb_dat_i[9]
  PIN wb_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 227.840 200.000 228.440 ;
    END
  END wb_dat_o[0]
  PIN wb_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 6.840 200.000 7.440 ;
    END
  END wb_dat_o[10]
  PIN wb_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 244.840 200.000 245.440 ;
    END
  END wb_dat_o[11]
  PIN wb_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 54.440 4.000 55.040 ;
    END
  END wb_dat_o[12]
  PIN wb_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 272.040 4.000 272.640 ;
    END
  END wb_dat_o[13]
  PIN wb_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 98.640 4.000 99.240 ;
    END
  END wb_dat_o[14]
  PIN wb_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END wb_dat_o[15]
  PIN wb_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 154.650 0.000 154.930 4.000 ;
    END
  END wb_dat_o[16]
  PIN wb_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 282.240 4.000 282.840 ;
    END
  END wb_dat_o[17]
  PIN wb_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.610 296.000 51.890 300.000 ;
    END
  END wb_dat_o[18]
  PIN wb_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.890 296.000 129.170 300.000 ;
    END
  END wb_dat_o[19]
  PIN wb_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 227.840 4.000 228.440 ;
    END
  END wb_dat_o[1]
  PIN wb_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 119.040 4.000 119.640 ;
    END
  END wb_dat_o[20]
  PIN wb_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.530 0.000 6.810 4.000 ;
    END
  END wb_dat_o[21]
  PIN wb_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.310 296.000 164.590 300.000 ;
    END
  END wb_dat_o[22]
  PIN wb_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.790 296.000 113.070 300.000 ;
    END
  END wb_dat_o[23]
  PIN wb_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.790 0.000 113.070 4.000 ;
    END
  END wb_dat_o[24]
  PIN wb_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.070 296.000 190.350 300.000 ;
    END
  END wb_dat_o[25]
  PIN wb_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 81.640 200.000 82.240 ;
    END
  END wb_dat_o[26]
  PIN wb_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 255.040 4.000 255.640 ;
    END
  END wb_dat_o[27]
  PIN wb_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 88.440 4.000 89.040 ;
    END
  END wb_dat_o[28]
  PIN wb_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.950 0.000 42.230 4.000 ;
    END
  END wb_dat_o[29]
  PIN wb_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.810 0.000 84.090 4.000 ;
    END
  END wb_dat_o[2]
  PIN wb_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.890 0.000 129.170 4.000 ;
    END
  END wb_dat_o[30]
  PIN wb_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 200.640 200.000 201.240 ;
    END
  END wb_dat_o[31]
  PIN wb_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.550 0.000 138.830 4.000 ;
    END
  END wb_dat_o[3]
  PIN wb_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.990 296.000 145.270 300.000 ;
    END
  END wb_dat_o[4]
  PIN wb_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.550 296.000 138.830 300.000 ;
    END
  END wb_dat_o[5]
  PIN wb_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 265.240 4.000 265.840 ;
    END
  END wb_dat_o[6]
  PIN wb_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 299.240 4.000 299.840 ;
    END
  END wb_dat_o[7]
  PIN wb_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.310 0.000 164.590 4.000 ;
    END
  END wb_dat_o[8]
  PIN wb_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 71.440 4.000 72.040 ;
    END
  END wb_dat_o[9]
  PIN wb_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 217.640 4.000 218.240 ;
    END
  END wb_stb_i
  PIN wb_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 163.240 200.000 163.840 ;
    END
  END wb_we_i
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 194.120 288.405 ;
      LAYER met1 ;
        RECT 0.070 10.640 199.940 289.980 ;
      LAYER met2 ;
        RECT 0.100 295.720 6.250 299.725 ;
        RECT 7.090 295.720 15.910 299.725 ;
        RECT 16.750 295.720 25.570 299.725 ;
        RECT 26.410 295.720 32.010 299.725 ;
        RECT 32.850 295.720 41.670 299.725 ;
        RECT 42.510 295.720 51.330 299.725 ;
        RECT 52.170 295.720 57.770 299.725 ;
        RECT 58.610 295.720 67.430 299.725 ;
        RECT 68.270 295.720 77.090 299.725 ;
        RECT 77.930 295.720 83.530 299.725 ;
        RECT 84.370 295.720 93.190 299.725 ;
        RECT 94.030 295.720 102.850 299.725 ;
        RECT 103.690 295.720 112.510 299.725 ;
        RECT 113.350 295.720 118.950 299.725 ;
        RECT 119.790 295.720 128.610 299.725 ;
        RECT 129.450 295.720 138.270 299.725 ;
        RECT 139.110 295.720 144.710 299.725 ;
        RECT 145.550 295.720 154.370 299.725 ;
        RECT 155.210 295.720 164.030 299.725 ;
        RECT 164.870 295.720 170.470 299.725 ;
        RECT 171.310 295.720 180.130 299.725 ;
        RECT 180.970 295.720 189.790 299.725 ;
        RECT 190.630 295.720 196.230 299.725 ;
        RECT 197.070 295.720 199.940 299.725 ;
        RECT 0.100 4.280 199.940 295.720 ;
        RECT 0.650 0.155 6.250 4.280 ;
        RECT 7.090 0.155 15.910 4.280 ;
        RECT 16.750 0.155 25.570 4.280 ;
        RECT 26.410 0.155 32.010 4.280 ;
        RECT 32.850 0.155 41.670 4.280 ;
        RECT 42.510 0.155 51.330 4.280 ;
        RECT 52.170 0.155 57.770 4.280 ;
        RECT 58.610 0.155 67.430 4.280 ;
        RECT 68.270 0.155 77.090 4.280 ;
        RECT 77.930 0.155 83.530 4.280 ;
        RECT 84.370 0.155 93.190 4.280 ;
        RECT 94.030 0.155 102.850 4.280 ;
        RECT 103.690 0.155 112.510 4.280 ;
        RECT 113.350 0.155 118.950 4.280 ;
        RECT 119.790 0.155 128.610 4.280 ;
        RECT 129.450 0.155 138.270 4.280 ;
        RECT 139.110 0.155 144.710 4.280 ;
        RECT 145.550 0.155 154.370 4.280 ;
        RECT 155.210 0.155 164.030 4.280 ;
        RECT 164.870 0.155 170.470 4.280 ;
        RECT 171.310 0.155 180.130 4.280 ;
        RECT 180.970 0.155 189.790 4.280 ;
        RECT 190.630 0.155 199.940 4.280 ;
      LAYER met3 ;
        RECT 4.400 298.840 199.575 299.705 ;
        RECT 4.000 293.440 199.575 298.840 ;
        RECT 4.400 292.040 195.600 293.440 ;
        RECT 4.000 283.240 199.575 292.040 ;
        RECT 4.400 281.840 195.600 283.240 ;
        RECT 4.000 273.040 199.575 281.840 ;
        RECT 4.400 271.640 195.600 273.040 ;
        RECT 4.000 266.240 199.575 271.640 ;
        RECT 4.400 264.840 195.600 266.240 ;
        RECT 4.000 256.040 199.575 264.840 ;
        RECT 4.400 254.640 195.600 256.040 ;
        RECT 4.000 245.840 199.575 254.640 ;
        RECT 4.400 244.440 195.600 245.840 ;
        RECT 4.000 239.040 199.575 244.440 ;
        RECT 4.400 237.640 195.600 239.040 ;
        RECT 4.000 228.840 199.575 237.640 ;
        RECT 4.400 227.440 195.600 228.840 ;
        RECT 4.000 218.640 199.575 227.440 ;
        RECT 4.400 217.240 195.600 218.640 ;
        RECT 4.000 211.840 199.575 217.240 ;
        RECT 4.400 210.440 195.600 211.840 ;
        RECT 4.000 201.640 199.575 210.440 ;
        RECT 4.400 200.240 195.600 201.640 ;
        RECT 4.000 191.440 199.575 200.240 ;
        RECT 4.400 190.040 195.600 191.440 ;
        RECT 4.000 181.240 199.575 190.040 ;
        RECT 4.400 179.840 195.600 181.240 ;
        RECT 4.000 174.440 199.575 179.840 ;
        RECT 4.400 173.040 195.600 174.440 ;
        RECT 4.000 164.240 199.575 173.040 ;
        RECT 4.400 162.840 195.600 164.240 ;
        RECT 4.000 154.040 199.575 162.840 ;
        RECT 4.400 152.640 195.600 154.040 ;
        RECT 4.000 147.240 199.575 152.640 ;
        RECT 4.400 145.840 195.600 147.240 ;
        RECT 4.000 137.040 199.575 145.840 ;
        RECT 4.400 135.640 195.600 137.040 ;
        RECT 4.000 126.840 199.575 135.640 ;
        RECT 4.400 125.440 195.600 126.840 ;
        RECT 4.000 120.040 199.575 125.440 ;
        RECT 4.400 118.640 195.600 120.040 ;
        RECT 4.000 109.840 199.575 118.640 ;
        RECT 4.400 108.440 195.600 109.840 ;
        RECT 4.000 99.640 199.575 108.440 ;
        RECT 4.400 98.240 195.600 99.640 ;
        RECT 4.000 89.440 199.575 98.240 ;
        RECT 4.400 88.040 195.600 89.440 ;
        RECT 4.000 82.640 199.575 88.040 ;
        RECT 4.400 81.240 195.600 82.640 ;
        RECT 4.000 72.440 199.575 81.240 ;
        RECT 4.400 71.040 195.600 72.440 ;
        RECT 4.000 62.240 199.575 71.040 ;
        RECT 4.400 60.840 195.600 62.240 ;
        RECT 4.000 55.440 199.575 60.840 ;
        RECT 4.400 54.040 195.600 55.440 ;
        RECT 4.000 45.240 199.575 54.040 ;
        RECT 4.400 43.840 195.600 45.240 ;
        RECT 4.000 35.040 199.575 43.840 ;
        RECT 4.400 33.640 195.600 35.040 ;
        RECT 4.000 28.240 199.575 33.640 ;
        RECT 4.400 26.840 195.600 28.240 ;
        RECT 4.000 18.040 199.575 26.840 ;
        RECT 4.400 16.640 195.600 18.040 ;
        RECT 4.000 7.840 199.575 16.640 ;
        RECT 4.400 6.440 195.600 7.840 ;
        RECT 4.000 1.040 199.575 6.440 ;
        RECT 4.000 0.175 195.600 1.040 ;
      LAYER met4 ;
        RECT 19.615 17.175 20.640 278.625 ;
        RECT 23.040 17.175 97.440 278.625 ;
        RECT 99.840 17.175 174.240 278.625 ;
        RECT 176.640 17.175 198.425 278.625 ;
  END
END trng_wb_wrapper
END LIBRARY

