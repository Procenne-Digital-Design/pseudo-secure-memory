VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_proj_example
  CLASS BLOCK ;
  FOREIGN user_proj_example ;
  ORIGIN 0.000 0.000 ;
  SIZE 1000.000 BY 1500.000 ;
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.930 1496.000 2.210 1500.000 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 115.090 1496.000 115.370 1500.000 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 126.130 1496.000 126.410 1500.000 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 137.630 1496.000 137.910 1500.000 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.670 1496.000 148.950 1500.000 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 160.170 1496.000 160.450 1500.000 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 171.670 1496.000 171.950 1500.000 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 182.710 1496.000 182.990 1500.000 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 194.210 1496.000 194.490 1500.000 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 205.710 1496.000 205.990 1500.000 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 216.750 1496.000 217.030 1500.000 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.970 1496.000 13.250 1500.000 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 228.250 1496.000 228.530 1500.000 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 239.290 1496.000 239.570 1500.000 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 250.790 1496.000 251.070 1500.000 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 262.290 1496.000 262.570 1500.000 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 273.330 1496.000 273.610 1500.000 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 284.830 1496.000 285.110 1500.000 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 295.870 1496.000 296.150 1500.000 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 307.370 1496.000 307.650 1500.000 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 318.870 1496.000 319.150 1500.000 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 329.910 1496.000 330.190 1500.000 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.470 1496.000 24.750 1500.000 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 341.410 1496.000 341.690 1500.000 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 352.450 1496.000 352.730 1500.000 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 363.950 1496.000 364.230 1500.000 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 375.450 1496.000 375.730 1500.000 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 386.490 1496.000 386.770 1500.000 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 397.990 1496.000 398.270 1500.000 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 409.490 1496.000 409.770 1500.000 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 420.530 1496.000 420.810 1500.000 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.510 1496.000 35.790 1500.000 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.010 1496.000 47.290 1500.000 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.510 1496.000 58.790 1500.000 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.550 1496.000 69.830 1500.000 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.050 1496.000 81.330 1500.000 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 92.090 1496.000 92.370 1500.000 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.590 1496.000 103.870 1500.000 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.610 1496.000 5.890 1500.000 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 118.770 1496.000 119.050 1500.000 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 129.810 1496.000 130.090 1500.000 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 141.310 1496.000 141.590 1500.000 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 152.810 1496.000 153.090 1500.000 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 163.850 1496.000 164.130 1500.000 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 175.350 1496.000 175.630 1500.000 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.390 1496.000 186.670 1500.000 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 197.890 1496.000 198.170 1500.000 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.390 1496.000 209.670 1500.000 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 220.430 1496.000 220.710 1500.000 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.650 1496.000 16.930 1500.000 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.930 1496.000 232.210 1500.000 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 243.430 1496.000 243.710 1500.000 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.470 1496.000 254.750 1500.000 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 265.970 1496.000 266.250 1500.000 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 277.010 1496.000 277.290 1500.000 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 288.510 1496.000 288.790 1500.000 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 300.010 1496.000 300.290 1500.000 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 311.050 1496.000 311.330 1500.000 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 322.550 1496.000 322.830 1500.000 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 333.590 1496.000 333.870 1500.000 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.150 1496.000 28.430 1500.000 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 345.090 1496.000 345.370 1500.000 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 356.590 1496.000 356.870 1500.000 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 367.630 1496.000 367.910 1500.000 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 379.130 1496.000 379.410 1500.000 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 390.170 1496.000 390.450 1500.000 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 401.670 1496.000 401.950 1500.000 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 413.170 1496.000 413.450 1500.000 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 424.210 1496.000 424.490 1500.000 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.650 1496.000 39.930 1500.000 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.690 1496.000 50.970 1500.000 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.190 1496.000 62.470 1500.000 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.230 1496.000 73.510 1500.000 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 84.730 1496.000 85.010 1500.000 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.230 1496.000 96.510 1500.000 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 107.270 1496.000 107.550 1500.000 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.290 1496.000 9.570 1500.000 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.450 1496.000 122.730 1500.000 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.950 1496.000 134.230 1500.000 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.990 1496.000 145.270 1500.000 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.490 1496.000 156.770 1500.000 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.530 1496.000 167.810 1500.000 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.030 1496.000 179.310 1500.000 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.530 1496.000 190.810 1500.000 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 201.570 1496.000 201.850 1500.000 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 213.070 1496.000 213.350 1500.000 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 224.570 1496.000 224.850 1500.000 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.790 1496.000 21.070 1500.000 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 235.610 1496.000 235.890 1500.000 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 247.110 1496.000 247.390 1500.000 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 258.150 1496.000 258.430 1500.000 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 269.650 1496.000 269.930 1500.000 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 281.150 1496.000 281.430 1500.000 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 292.190 1496.000 292.470 1500.000 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 303.690 1496.000 303.970 1500.000 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 314.730 1496.000 315.010 1500.000 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 326.230 1496.000 326.510 1500.000 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 337.730 1496.000 338.010 1500.000 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.830 1496.000 32.110 1500.000 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 348.770 1496.000 349.050 1500.000 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 360.270 1496.000 360.550 1500.000 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 371.310 1496.000 371.590 1500.000 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 382.810 1496.000 383.090 1500.000 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 394.310 1496.000 394.590 1500.000 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 405.350 1496.000 405.630 1500.000 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 416.850 1496.000 417.130 1500.000 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 428.350 1496.000 428.630 1500.000 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.330 1496.000 43.610 1500.000 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.370 1496.000 54.650 1500.000 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.870 1496.000 66.150 1500.000 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.370 1496.000 77.650 1500.000 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.410 1496.000 88.690 1500.000 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.910 1496.000 100.190 1500.000 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.950 1496.000 111.230 1500.000 ;
    END
  END io_out[9]
  PIN irq[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 395.690 0.000 395.970 4.000 ;
    END
  END irq[0]
  PIN irq[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 399.370 0.000 399.650 4.000 ;
    END
  END irq[1]
  PIN irq[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 403.050 0.000 403.330 4.000 ;
    END
  END irq[2]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 18.400 4.000 19.000 ;
    END
  END la_data_in[0]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 903.530 1496.000 903.810 1500.000 ;
    END
  END la_data_in[100]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 915.030 1496.000 915.310 1500.000 ;
    END
  END la_data_in[101]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 1296.120 1000.000 1296.720 ;
    END
  END la_data_in[102]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 922.390 1496.000 922.670 1500.000 ;
    END
  END la_data_in[103]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 1315.840 1000.000 1316.440 ;
    END
  END la_data_in[104]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 920.090 0.000 920.370 4.000 ;
    END
  END la_data_in[105]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 930.210 1496.000 930.490 1500.000 ;
    END
  END la_data_in[106]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 1335.560 1000.000 1336.160 ;
    END
  END la_data_in[107]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 933.890 1496.000 934.170 1500.000 ;
    END
  END la_data_in[108]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 1355.280 1000.000 1355.880 ;
    END
  END la_data_in[109]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 536.910 0.000 537.190 4.000 ;
    END
  END la_data_in[10]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 941.250 1496.000 941.530 1500.000 ;
    END
  END la_data_in[110]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 949.530 0.000 949.810 4.000 ;
    END
  END la_data_in[111]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 1375.680 1000.000 1376.280 ;
    END
  END la_data_in[112]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 949.070 1496.000 949.350 1500.000 ;
    END
  END la_data_in[113]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 961.030 0.000 961.310 4.000 ;
    END
  END la_data_in[114]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 956.430 1496.000 956.710 1500.000 ;
    END
  END la_data_in[115]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 964.710 0.000 964.990 4.000 ;
    END
  END la_data_in[116]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 968.390 0.000 968.670 4.000 ;
    END
  END la_data_in[117]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 971.610 1496.000 971.890 1500.000 ;
    END
  END la_data_in[118]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 979.430 0.000 979.710 4.000 ;
    END
  END la_data_in[119]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 330.520 4.000 331.120 ;
    END
  END la_data_in[11]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1418.520 4.000 1419.120 ;
    END
  END la_data_in[120]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1443.680 4.000 1444.280 ;
    END
  END la_data_in[121]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 1454.560 1000.000 1455.160 ;
    END
  END la_data_in[122]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 1474.960 1000.000 1475.560 ;
    END
  END la_data_in[123]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 986.790 1496.000 987.070 1500.000 ;
    END
  END la_data_in[124]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 1494.680 1000.000 1495.280 ;
    END
  END la_data_in[125]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 994.150 0.000 994.430 4.000 ;
    END
  END la_data_in[126]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 997.830 1496.000 998.110 1500.000 ;
    END
  END la_data_in[127]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 343.440 4.000 344.040 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 556.230 1496.000 556.510 1500.000 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 355.680 4.000 356.280 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 582.910 1496.000 583.190 1500.000 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 600.390 0.000 600.670 4.000 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 431.840 1000.000 432.440 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 418.240 4.000 418.840 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 481.480 1000.000 482.080 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 421.910 0.000 422.190 4.000 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 501.200 1000.000 501.800 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 493.040 4.000 493.640 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 639.490 1496.000 639.770 1500.000 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 656.050 0.000 656.330 4.000 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 570.560 1000.000 571.160 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 543.360 4.000 543.960 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 669.850 1496.000 670.130 1500.000 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 580.760 4.000 581.360 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 605.920 4.000 606.520 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 690.240 1000.000 690.840 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 436.630 0.000 436.910 4.000 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 699.750 1496.000 700.030 1500.000 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 749.400 1000.000 750.000 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 719.070 0.000 719.350 4.000 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 726.430 0.000 726.710 4.000 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 769.120 1000.000 769.720 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 741.610 0.000 741.890 4.000 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 722.290 1496.000 722.570 1500.000 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 768.440 4.000 769.040 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 779.320 1000.000 779.920 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 789.520 1000.000 790.120 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 451.350 0.000 451.630 4.000 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 730.110 1496.000 730.390 1500.000 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 805.840 4.000 806.440 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 763.690 0.000 763.970 4.000 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 745.290 1496.000 745.570 1500.000 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 771.050 0.000 771.330 4.000 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 778.870 0.000 779.150 4.000 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 843.240 4.000 843.840 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 856.160 4.000 856.760 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 880.640 4.000 881.240 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 828.960 1000.000 829.560 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 130.600 4.000 131.200 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 756.330 1496.000 756.610 1500.000 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 760.010 1496.000 760.290 1500.000 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 905.800 4.000 906.400 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 930.960 4.000 931.560 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 767.830 1496.000 768.110 1500.000 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 888.800 1000.000 889.400 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 908.520 1000.000 909.120 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 928.240 1000.000 928.840 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 947.960 1000.000 948.560 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 958.160 1000.000 958.760 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 480.790 1496.000 481.070 1500.000 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 815.670 0.000 815.950 4.000 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 988.080 1000.000 988.680 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 783.010 1496.000 783.290 1500.000 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1018.680 4.000 1019.280 ;
    END
  END la_data_in[63]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 827.170 0.000 827.450 4.000 ;
    END
  END la_data_in[64]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 790.370 1496.000 790.650 1500.000 ;
    END
  END la_data_in[65]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 797.730 1496.000 798.010 1500.000 ;
    END
  END la_data_in[66]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1043.160 4.000 1043.760 ;
    END
  END la_data_in[67]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1056.080 4.000 1056.680 ;
    END
  END la_data_in[68]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 1037.720 1000.000 1038.320 ;
    END
  END la_data_in[69]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 242.800 1000.000 243.400 ;
    END
  END la_data_in[6]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 841.890 0.000 842.170 4.000 ;
    END
  END la_data_in[70]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 1047.240 1000.000 1047.840 ;
    END
  END la_data_in[71]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 845.570 0.000 845.850 4.000 ;
    END
  END la_data_in[72]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1105.720 4.000 1106.320 ;
    END
  END la_data_in[73]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 1067.640 1000.000 1068.240 ;
    END
  END la_data_in[74]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1118.640 4.000 1119.240 ;
    END
  END la_data_in[75]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 1087.360 1000.000 1087.960 ;
    END
  END la_data_in[76]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 1097.560 1000.000 1098.160 ;
    END
  END la_data_in[77]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 863.970 0.000 864.250 4.000 ;
    END
  END la_data_in[78]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 835.910 1496.000 836.190 1500.000 ;
    END
  END la_data_in[79]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 495.970 0.000 496.250 4.000 ;
    END
  END la_data_in[7]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1168.280 4.000 1168.880 ;
    END
  END la_data_in[80]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 839.590 1496.000 839.870 1500.000 ;
    END
  END la_data_in[81]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 843.270 1496.000 843.550 1500.000 ;
    END
  END la_data_in[82]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 1126.800 1000.000 1127.400 ;
    END
  END la_data_in[83]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 882.830 0.000 883.110 4.000 ;
    END
  END la_data_in[84]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 858.450 1496.000 858.730 1500.000 ;
    END
  END la_data_in[85]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 1147.200 1000.000 1147.800 ;
    END
  END la_data_in[86]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 886.510 0.000 886.790 4.000 ;
    END
  END la_data_in[87]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 1166.920 1000.000 1167.520 ;
    END
  END la_data_in[88]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 1176.440 1000.000 1177.040 ;
    END
  END la_data_in[89]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 511.150 0.000 511.430 4.000 ;
    END
  END la_data_in[8]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 877.310 1496.000 877.590 1500.000 ;
    END
  END la_data_in[90]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 1196.840 1000.000 1197.440 ;
    END
  END la_data_in[91]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 1226.080 1000.000 1226.680 ;
    END
  END la_data_in[92]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 1236.280 1000.000 1236.880 ;
    END
  END la_data_in[93]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 888.350 1496.000 888.630 1500.000 ;
    END
  END la_data_in[94]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1268.240 4.000 1268.840 ;
    END
  END la_data_in[95]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 896.170 1496.000 896.450 1500.000 ;
    END
  END la_data_in[96]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 1266.200 1000.000 1266.800 ;
    END
  END la_data_in[97]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 1275.720 1000.000 1276.320 ;
    END
  END la_data_in[98]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1318.560 4.000 1319.160 ;
    END
  END la_data_in[99]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 499.650 1496.000 499.930 1500.000 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 414.550 0.000 414.830 4.000 ;
    END
  END la_data_out[0]
  PIN la_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 907.210 1496.000 907.490 1500.000 ;
    END
  END la_data_out[100]
  PIN la_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1330.800 4.000 1331.400 ;
    END
  END la_data_out[101]
  PIN la_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 916.410 0.000 916.690 4.000 ;
    END
  END la_data_out[102]
  PIN la_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1343.720 4.000 1344.320 ;
    END
  END la_data_out[103]
  PIN la_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1368.200 4.000 1368.800 ;
    END
  END la_data_out[104]
  PIN la_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 1326.040 1000.000 1326.640 ;
    END
  END la_data_out[105]
  PIN la_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 927.450 0.000 927.730 4.000 ;
    END
  END la_data_out[106]
  PIN la_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 931.130 0.000 931.410 4.000 ;
    END
  END la_data_out[107]
  PIN la_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 934.810 0.000 935.090 4.000 ;
    END
  END la_data_out[108]
  PIN la_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 942.170 0.000 942.450 4.000 ;
    END
  END la_data_out[109]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 514.830 1496.000 515.110 1500.000 ;
    END
  END la_data_out[10]
  PIN la_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 945.850 0.000 946.130 4.000 ;
    END
  END la_data_out[110]
  PIN la_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1393.360 4.000 1393.960 ;
    END
  END la_data_out[111]
  PIN la_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 953.210 0.000 953.490 4.000 ;
    END
  END la_data_out[112]
  PIN la_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 957.350 0.000 957.630 4.000 ;
    END
  END la_data_out[113]
  PIN la_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 1395.400 1000.000 1396.000 ;
    END
  END la_data_out[114]
  PIN la_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 1415.120 1000.000 1415.720 ;
    END
  END la_data_out[115]
  PIN la_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 963.790 1496.000 964.070 1500.000 ;
    END
  END la_data_out[116]
  PIN la_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 967.930 1496.000 968.210 1500.000 ;
    END
  END la_data_out[117]
  PIN la_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 975.750 0.000 976.030 4.000 ;
    END
  END la_data_out[118]
  PIN la_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 975.290 1496.000 975.570 1500.000 ;
    END
  END la_data_out[119]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 526.330 1496.000 526.610 1500.000 ;
    END
  END la_data_out[11]
  PIN la_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1430.760 4.000 1431.360 ;
    END
  END la_data_out[120]
  PIN la_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 978.970 1496.000 979.250 1500.000 ;
    END
  END la_data_out[121]
  PIN la_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 1464.760 1000.000 1465.360 ;
    END
  END la_data_out[122]
  PIN la_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1468.160 4.000 1468.760 ;
    END
  END la_data_out[123]
  PIN la_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 1484.480 1000.000 1485.080 ;
    END
  END la_data_out[124]
  PIN la_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 986.790 0.000 987.070 4.000 ;
    END
  END la_data_out[125]
  PIN la_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 994.150 1496.000 994.430 1500.000 ;
    END
  END la_data_out[126]
  PIN la_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1481.080 4.000 1481.680 ;
    END
  END la_data_out[127]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 541.510 1496.000 541.790 1500.000 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 570.490 0.000 570.770 4.000 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 571.410 1496.000 571.690 1500.000 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 401.920 1000.000 402.520 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 380.840 4.000 381.440 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 604.070 0.000 604.350 4.000 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 431.160 4.000 431.760 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 615.110 0.000 615.390 4.000 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 34.040 1000.000 34.640 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 626.150 0.000 626.430 4.000 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 511.400 1000.000 512.000 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 520.920 1000.000 521.520 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 518.200 4.000 518.800 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 670.770 0.000 671.050 4.000 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 610.680 1000.000 611.280 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 630.400 1000.000 631.000 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 650.120 1000.000 650.720 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 618.160 4.000 618.760 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 699.760 1000.000 700.360 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 440.310 0.000 440.590 4.000 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 729.680 1000.000 730.280 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 711.250 1496.000 711.530 1500.000 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 722.750 0.000 723.030 4.000 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 730.570 0.000 730.850 4.000 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 734.250 0.000 734.530 4.000 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 731.040 4.000 731.640 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 743.280 4.000 743.880 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 748.970 0.000 749.250 4.000 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 752.650 0.000 752.930 4.000 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 726.430 1496.000 726.710 1500.000 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 133.320 1000.000 133.920 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 733.790 1496.000 734.070 1500.000 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 737.470 1496.000 737.750 1500.000 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 741.150 1496.000 741.430 1500.000 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 799.040 1000.000 799.640 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 775.190 0.000 775.470 4.000 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 782.550 0.000 782.830 4.000 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 786.230 0.000 786.510 4.000 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 818.760 1000.000 819.360 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 793.590 0.000 793.870 4.000 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 839.160 1000.000 839.760 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 466.530 0.000 466.810 4.000 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 848.680 1000.000 849.280 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 764.150 1496.000 764.430 1500.000 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 858.880 1000.000 859.480 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 943.200 4.000 943.800 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 878.600 1000.000 879.200 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 804.630 0.000 804.910 4.000 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 918.720 1000.000 919.320 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 956.120 4.000 956.720 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 811.990 0.000 812.270 4.000 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 968.360 1000.000 968.960 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 206.080 4.000 206.680 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 778.870 1496.000 779.150 1500.000 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 819.350 0.000 819.630 4.000 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 993.520 4.000 994.120 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 823.490 0.000 823.770 4.000 ;
    END
  END la_data_out[63]
  PIN la_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 997.600 1000.000 998.200 ;
    END
  END la_data_out[64]
  PIN la_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 794.050 1496.000 794.330 1500.000 ;
    END
  END la_data_out[65]
  PIN la_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 801.870 1496.000 802.150 1500.000 ;
    END
  END la_data_out[66]
  PIN la_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 834.530 0.000 834.810 4.000 ;
    END
  END la_data_out[67]
  PIN la_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 1027.520 1000.000 1028.120 ;
    END
  END la_data_out[68]
  PIN la_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1080.560 4.000 1081.160 ;
    END
  END la_data_out[69]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 253.000 1000.000 253.600 ;
    END
  END la_data_out[6]
  PIN la_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 805.550 1496.000 805.830 1500.000 ;
    END
  END la_data_out[70]
  PIN la_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 812.910 1496.000 813.190 1500.000 ;
    END
  END la_data_out[71]
  PIN la_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1093.480 4.000 1094.080 ;
    END
  END la_data_out[72]
  PIN la_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 852.930 0.000 853.210 4.000 ;
    END
  END la_data_out[73]
  PIN la_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 856.610 0.000 856.890 4.000 ;
    END
  END la_data_out[74]
  PIN la_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 824.410 1496.000 824.690 1500.000 ;
    END
  END la_data_out[75]
  PIN la_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1130.880 4.000 1131.480 ;
    END
  END la_data_out[76]
  PIN la_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 828.090 1496.000 828.370 1500.000 ;
    END
  END la_data_out[77]
  PIN la_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 831.770 1496.000 832.050 1500.000 ;
    END
  END la_data_out[78]
  PIN la_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1156.040 4.000 1156.640 ;
    END
  END la_data_out[79]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 272.720 1000.000 273.320 ;
    END
  END la_data_out[7]
  PIN la_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1181.200 4.000 1181.800 ;
    END
  END la_data_out[80]
  PIN la_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 871.790 0.000 872.070 4.000 ;
    END
  END la_data_out[81]
  PIN la_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 846.950 1496.000 847.230 1500.000 ;
    END
  END la_data_out[82]
  PIN la_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 879.150 0.000 879.430 4.000 ;
    END
  END la_data_out[83]
  PIN la_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1193.440 4.000 1194.040 ;
    END
  END la_data_out[84]
  PIN la_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1205.680 4.000 1206.280 ;
    END
  END la_data_out[85]
  PIN la_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 865.810 1496.000 866.090 1500.000 ;
    END
  END la_data_out[86]
  PIN la_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 869.490 1496.000 869.770 1500.000 ;
    END
  END la_data_out[87]
  PIN la_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1218.600 4.000 1219.200 ;
    END
  END la_data_out[88]
  PIN la_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 1186.640 1000.000 1187.240 ;
    END
  END la_data_out[89]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 302.640 1000.000 303.240 ;
    END
  END la_data_out[8]
  PIN la_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 880.990 1496.000 881.270 1500.000 ;
    END
  END la_data_out[90]
  PIN la_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 1206.360 1000.000 1206.960 ;
    END
  END la_data_out[91]
  PIN la_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1243.080 4.000 1243.680 ;
    END
  END la_data_out[92]
  PIN la_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 884.670 1496.000 884.950 1500.000 ;
    END
  END la_data_out[93]
  PIN la_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 892.490 1496.000 892.770 1500.000 ;
    END
  END la_data_out[94]
  PIN la_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 897.550 0.000 897.830 4.000 ;
    END
  END la_data_out[95]
  PIN la_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 899.850 1496.000 900.130 1500.000 ;
    END
  END la_data_out[96]
  PIN la_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1293.400 4.000 1294.000 ;
    END
  END la_data_out[97]
  PIN la_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 908.590 0.000 908.870 4.000 ;
    END
  END la_data_out[98]
  PIN la_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 912.730 0.000 913.010 4.000 ;
    END
  END la_data_out[99]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 529.550 0.000 529.830 4.000 ;
    END
  END la_data_out[9]
  PIN la_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 4.800 1000.000 5.400 ;
    END
  END la_oenb[0]
  PIN la_oenb[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 911.350 1496.000 911.630 1500.000 ;
    END
  END la_oenb[100]
  PIN la_oenb[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 918.710 1496.000 918.990 1500.000 ;
    END
  END la_oenb[101]
  PIN la_oenb[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 1305.640 1000.000 1306.240 ;
    END
  END la_oenb[102]
  PIN la_oenb[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1355.960 4.000 1356.560 ;
    END
  END la_oenb[103]
  PIN la_oenb[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 926.070 1496.000 926.350 1500.000 ;
    END
  END la_oenb[104]
  PIN la_oenb[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 923.770 0.000 924.050 4.000 ;
    END
  END la_oenb[105]
  PIN la_oenb[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1381.120 4.000 1381.720 ;
    END
  END la_oenb[106]
  PIN la_oenb[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 1345.760 1000.000 1346.360 ;
    END
  END la_oenb[107]
  PIN la_oenb[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 938.490 0.000 938.770 4.000 ;
    END
  END la_oenb[108]
  PIN la_oenb[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 937.570 1496.000 937.850 1500.000 ;
    END
  END la_oenb[109]
  PIN la_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 540.590 0.000 540.870 4.000 ;
    END
  END la_oenb[10]
  PIN la_oenb[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 1365.480 1000.000 1366.080 ;
    END
  END la_oenb[110]
  PIN la_oenb[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 944.930 1496.000 945.210 1500.000 ;
    END
  END la_oenb[111]
  PIN la_oenb[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 1385.200 1000.000 1385.800 ;
    END
  END la_oenb[112]
  PIN la_oenb[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 952.750 1496.000 953.030 1500.000 ;
    END
  END la_oenb[113]
  PIN la_oenb[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 1404.920 1000.000 1405.520 ;
    END
  END la_oenb[114]
  PIN la_oenb[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 960.110 1496.000 960.390 1500.000 ;
    END
  END la_oenb[115]
  PIN la_oenb[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 1425.320 1000.000 1425.920 ;
    END
  END la_oenb[116]
  PIN la_oenb[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 972.070 0.000 972.350 4.000 ;
    END
  END la_oenb[117]
  PIN la_oenb[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 1434.840 1000.000 1435.440 ;
    END
  END la_oenb[118]
  PIN la_oenb[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1405.600 4.000 1406.200 ;
    END
  END la_oenb[119]
  PIN la_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 530.010 1496.000 530.290 1500.000 ;
    END
  END la_oenb[11]
  PIN la_oenb[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 1445.040 1000.000 1445.640 ;
    END
  END la_oenb[120]
  PIN la_oenb[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 983.110 0.000 983.390 4.000 ;
    END
  END la_oenb[121]
  PIN la_oenb[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1455.920 4.000 1456.520 ;
    END
  END la_oenb[122]
  PIN la_oenb[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 982.650 1496.000 982.930 1500.000 ;
    END
  END la_oenb[123]
  PIN la_oenb[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 990.470 1496.000 990.750 1500.000 ;
    END
  END la_oenb[124]
  PIN la_oenb[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 990.470 0.000 990.750 4.000 ;
    END
  END la_oenb[125]
  PIN la_oenb[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 997.830 0.000 998.110 4.000 ;
    END
  END la_oenb[126]
  PIN la_oenb[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1493.320 4.000 1493.920 ;
    END
  END la_oenb[127]
  PIN la_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 559.450 0.000 559.730 4.000 ;
    END
  END la_oenb[12]
  PIN la_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 560.370 1496.000 560.650 1500.000 ;
    END
  END la_oenb[13]
  PIN la_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 575.090 1496.000 575.370 1500.000 ;
    END
  END la_oenb[14]
  PIN la_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 588.890 0.000 589.170 4.000 ;
    END
  END la_oenb[15]
  PIN la_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 590.270 1496.000 590.550 1500.000 ;
    END
  END la_oenb[16]
  PIN la_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 441.360 1000.000 441.960 ;
    END
  END la_oenb[17]
  PIN la_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 607.750 0.000 608.030 4.000 ;
    END
  END la_oenb[18]
  PIN la_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 618.790 0.000 619.070 4.000 ;
    END
  END la_oenb[19]
  PIN la_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 425.590 0.000 425.870 4.000 ;
    END
  END la_oenb[1]
  PIN la_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 624.310 1496.000 624.590 1500.000 ;
    END
  END la_oenb[20]
  PIN la_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 627.990 1496.000 628.270 1500.000 ;
    END
  END la_oenb[21]
  PIN la_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 652.370 0.000 652.650 4.000 ;
    END
  END la_oenb[22]
  PIN la_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 659.730 0.000 660.010 4.000 ;
    END
  END la_oenb[23]
  PIN la_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 654.670 1496.000 654.950 1500.000 ;
    END
  END la_oenb[24]
  PIN la_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 620.200 1000.000 620.800 ;
    END
  END la_oenb[25]
  PIN la_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 639.920 1000.000 640.520 ;
    END
  END la_oenb[26]
  PIN la_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 593.680 4.000 594.280 ;
    END
  END la_oenb[27]
  PIN la_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 688.710 1496.000 688.990 1500.000 ;
    END
  END la_oenb[28]
  PIN la_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 709.960 1000.000 710.560 ;
    END
  END la_oenb[29]
  PIN la_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 93.200 4.000 93.800 ;
    END
  END la_oenb[2]
  PIN la_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 703.430 1496.000 703.710 1500.000 ;
    END
  END la_oenb[30]
  PIN la_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 714.930 1496.000 715.210 1500.000 ;
    END
  END la_oenb[31]
  PIN la_oenb[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 718.120 4.000 718.720 ;
    END
  END la_oenb[32]
  PIN la_oenb[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 718.610 1496.000 718.890 1500.000 ;
    END
  END la_oenb[33]
  PIN la_oenb[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 737.930 0.000 738.210 4.000 ;
    END
  END la_oenb[34]
  PIN la_oenb[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 745.290 0.000 745.570 4.000 ;
    END
  END la_oenb[35]
  PIN la_oenb[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 756.200 4.000 756.800 ;
    END
  END la_oenb[36]
  PIN la_oenb[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 780.680 4.000 781.280 ;
    END
  END la_oenb[37]
  PIN la_oenb[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 756.330 0.000 756.610 4.000 ;
    END
  END la_oenb[38]
  PIN la_oenb[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 793.600 4.000 794.200 ;
    END
  END la_oenb[39]
  PIN la_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 466.070 1496.000 466.350 1500.000 ;
    END
  END la_oenb[3]
  PIN la_oenb[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 760.010 0.000 760.290 4.000 ;
    END
  END la_oenb[40]
  PIN la_oenb[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 818.080 4.000 818.680 ;
    END
  END la_oenb[41]
  PIN la_oenb[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 767.370 0.000 767.650 4.000 ;
    END
  END la_oenb[42]
  PIN la_oenb[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 809.240 1000.000 809.840 ;
    END
  END la_oenb[43]
  PIN la_oenb[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 831.000 4.000 831.600 ;
    END
  END la_oenb[44]
  PIN la_oenb[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 748.970 1496.000 749.250 1500.000 ;
    END
  END la_oenb[45]
  PIN la_oenb[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 789.910 0.000 790.190 4.000 ;
    END
  END la_oenb[46]
  PIN la_oenb[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 868.400 4.000 869.000 ;
    END
  END la_oenb[47]
  PIN la_oenb[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 893.560 4.000 894.160 ;
    END
  END la_oenb[48]
  PIN la_oenb[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 752.650 1496.000 752.930 1500.000 ;
    END
  END la_oenb[49]
  PIN la_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 477.110 1496.000 477.390 1500.000 ;
    END
  END la_oenb[4]
  PIN la_oenb[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 797.270 0.000 797.550 4.000 ;
    END
  END la_oenb[50]
  PIN la_oenb[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 800.950 0.000 801.230 4.000 ;
    END
  END la_oenb[51]
  PIN la_oenb[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 918.040 4.000 918.640 ;
    END
  END la_oenb[52]
  PIN la_oenb[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 869.080 1000.000 869.680 ;
    END
  END la_oenb[53]
  PIN la_oenb[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 771.510 1496.000 771.790 1500.000 ;
    END
  END la_oenb[54]
  PIN la_oenb[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 898.320 1000.000 898.920 ;
    END
  END la_oenb[55]
  PIN la_oenb[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 808.310 0.000 808.590 4.000 ;
    END
  END la_oenb[56]
  PIN la_oenb[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 938.440 1000.000 939.040 ;
    END
  END la_oenb[57]
  PIN la_oenb[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 775.190 1496.000 775.470 1500.000 ;
    END
  END la_oenb[58]
  PIN la_oenb[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 977.880 1000.000 978.480 ;
    END
  END la_oenb[59]
  PIN la_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 193.160 1000.000 193.760 ;
    END
  END la_oenb[5]
  PIN la_oenb[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 968.360 4.000 968.960 ;
    END
  END la_oenb[60]
  PIN la_oenb[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 980.600 4.000 981.200 ;
    END
  END la_oenb[61]
  PIN la_oenb[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1005.760 4.000 1006.360 ;
    END
  END la_oenb[62]
  PIN la_oenb[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 786.690 1496.000 786.970 1500.000 ;
    END
  END la_oenb[63]
  PIN la_oenb[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1030.920 4.000 1031.520 ;
    END
  END la_oenb[64]
  PIN la_oenb[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 830.850 0.000 831.130 4.000 ;
    END
  END la_oenb[65]
  PIN la_oenb[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 1007.800 1000.000 1008.400 ;
    END
  END la_oenb[66]
  PIN la_oenb[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 1018.000 1000.000 1018.600 ;
    END
  END la_oenb[67]
  PIN la_oenb[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1068.320 4.000 1068.920 ;
    END
  END la_oenb[68]
  PIN la_oenb[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 838.210 0.000 838.490 4.000 ;
    END
  END la_oenb[69]
  PIN la_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 230.560 4.000 231.160 ;
    END
  END la_oenb[6]
  PIN la_oenb[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 809.230 1496.000 809.510 1500.000 ;
    END
  END la_oenb[70]
  PIN la_oenb[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 1057.440 1000.000 1058.040 ;
    END
  END la_oenb[71]
  PIN la_oenb[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 849.250 0.000 849.530 4.000 ;
    END
  END la_oenb[72]
  PIN la_oenb[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 817.050 1496.000 817.330 1500.000 ;
    END
  END la_oenb[73]
  PIN la_oenb[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 820.730 1496.000 821.010 1500.000 ;
    END
  END la_oenb[74]
  PIN la_oenb[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 1077.160 1000.000 1077.760 ;
    END
  END la_oenb[75]
  PIN la_oenb[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1143.120 4.000 1143.720 ;
    END
  END la_oenb[76]
  PIN la_oenb[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 860.290 0.000 860.570 4.000 ;
    END
  END la_oenb[77]
  PIN la_oenb[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 1107.080 1000.000 1107.680 ;
    END
  END la_oenb[78]
  PIN la_oenb[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 868.110 0.000 868.390 4.000 ;
    END
  END la_oenb[79]
  PIN la_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 268.640 4.000 269.240 ;
    END
  END la_oenb[7]
  PIN la_oenb[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 1117.280 1000.000 1117.880 ;
    END
  END la_oenb[80]
  PIN la_oenb[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 875.470 0.000 875.750 4.000 ;
    END
  END la_oenb[81]
  PIN la_oenb[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 850.630 1496.000 850.910 1500.000 ;
    END
  END la_oenb[82]
  PIN la_oenb[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 854.770 1496.000 855.050 1500.000 ;
    END
  END la_oenb[83]
  PIN la_oenb[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 1137.000 1000.000 1137.600 ;
    END
  END la_oenb[84]
  PIN la_oenb[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 862.130 1496.000 862.410 1500.000 ;
    END
  END la_oenb[85]
  PIN la_oenb[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 1156.720 1000.000 1157.320 ;
    END
  END la_oenb[86]
  PIN la_oenb[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 873.630 1496.000 873.910 1500.000 ;
    END
  END la_oenb[87]
  PIN la_oenb[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1230.840 4.000 1231.440 ;
    END
  END la_oenb[88]
  PIN la_oenb[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 890.190 0.000 890.470 4.000 ;
    END
  END la_oenb[89]
  PIN la_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 495.970 1496.000 496.250 1500.000 ;
    END
  END la_oenb[8]
  PIN la_oenb[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 893.870 0.000 894.150 4.000 ;
    END
  END la_oenb[90]
  PIN la_oenb[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 1216.560 1000.000 1217.160 ;
    END
  END la_oenb[91]
  PIN la_oenb[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1256.000 4.000 1256.600 ;
    END
  END la_oenb[92]
  PIN la_oenb[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 1246.480 1000.000 1247.080 ;
    END
  END la_oenb[93]
  PIN la_oenb[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 1256.000 1000.000 1256.600 ;
    END
  END la_oenb[94]
  PIN la_oenb[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 901.230 0.000 901.510 4.000 ;
    END
  END la_oenb[95]
  PIN la_oenb[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1281.160 4.000 1281.760 ;
    END
  END la_oenb[96]
  PIN la_oenb[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 904.910 0.000 905.190 4.000 ;
    END
  END la_oenb[97]
  PIN la_oenb[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1305.640 4.000 1306.240 ;
    END
  END la_oenb[98]
  PIN la_oenb[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 1285.920 1000.000 1286.520 ;
    END
  END la_oenb[99]
  PIN la_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 533.230 0.000 533.510 4.000 ;
    END
  END la_oenb[9]
  PIN sram_addr_a[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 14.320 1000.000 14.920 ;
    END
  END sram_addr_a[0]
  PIN sram_addr_a[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 80.960 4.000 81.560 ;
    END
  END sram_addr_a[1]
  PIN sram_addr_a[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 458.250 1496.000 458.530 1500.000 ;
    END
  END sram_addr_a[2]
  PIN sram_addr_a[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 455.030 0.000 455.310 4.000 ;
    END
  END sram_addr_a[3]
  PIN sram_addr_a[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 143.520 4.000 144.120 ;
    END
  END sram_addr_a[4]
  PIN sram_addr_a[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 473.890 0.000 474.170 4.000 ;
    END
  END sram_addr_a[5]
  PIN sram_addr_a[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 262.520 1000.000 263.120 ;
    END
  END sram_addr_a[6]
  PIN sram_addr_a[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 499.650 0.000 499.930 4.000 ;
    END
  END sram_addr_a[7]
  PIN sram_addr_a[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 306.040 4.000 306.640 ;
    END
  END sram_addr_a[8]
  PIN sram_addr_b[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 30.640 4.000 31.240 ;
    END
  END sram_addr_b[0]
  PIN sram_addr_b[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 44.240 1000.000 44.840 ;
    END
  END sram_addr_b[1]
  PIN sram_addr_b[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 93.880 1000.000 94.480 ;
    END
  END sram_addr_b[2]
  PIN sram_addr_b[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 143.520 1000.000 144.120 ;
    END
  END sram_addr_b[3]
  PIN sram_addr_b[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 155.760 4.000 156.360 ;
    END
  END sram_addr_b[4]
  PIN sram_addr_b[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 203.360 1000.000 203.960 ;
    END
  END sram_addr_b[5]
  PIN sram_addr_b[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 243.480 4.000 244.080 ;
    END
  END sram_addr_b[6]
  PIN sram_addr_b[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 492.290 1496.000 492.570 1500.000 ;
    END
  END sram_addr_b[7]
  PIN sram_addr_b[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 514.830 0.000 515.110 4.000 ;
    END
  END sram_addr_b[8]
  PIN sram_csb_a
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 6.160 4.000 6.760 ;
    END
  END sram_csb_a
  PIN sram_csb_b
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 406.730 0.000 407.010 4.000 ;
    END
  END sram_csb_b
  PIN sram_din_b[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 43.560 4.000 44.160 ;
    END
  END sram_din_b[0]
  PIN sram_din_b[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 318.280 4.000 318.880 ;
    END
  END sram_din_b[10]
  PIN sram_din_b[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 533.690 1496.000 533.970 1500.000 ;
    END
  END sram_din_b[11]
  PIN sram_din_b[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 563.130 0.000 563.410 4.000 ;
    END
  END sram_din_b[12]
  PIN sram_din_b[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 564.050 1496.000 564.330 1500.000 ;
    END
  END sram_din_b[13]
  PIN sram_din_b[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 577.850 0.000 578.130 4.000 ;
    END
  END sram_din_b[14]
  PIN sram_din_b[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 368.600 4.000 369.200 ;
    END
  END sram_din_b[15]
  PIN sram_din_b[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 393.080 4.000 393.680 ;
    END
  END sram_din_b[16]
  PIN sram_din_b[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 451.560 1000.000 452.160 ;
    END
  END sram_din_b[17]
  PIN sram_din_b[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 609.130 1496.000 609.410 1500.000 ;
    END
  END sram_din_b[18]
  PIN sram_din_b[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 622.470 0.000 622.750 4.000 ;
    END
  END sram_din_b[19]
  PIN sram_din_b[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 429.270 0.000 429.550 4.000 ;
    END
  END sram_din_b[1]
  PIN sram_din_b[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 629.830 0.000 630.110 4.000 ;
    END
  END sram_din_b[20]
  PIN sram_din_b[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 645.010 0.000 645.290 4.000 ;
    END
  END sram_din_b[21]
  PIN sram_din_b[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 531.120 1000.000 531.720 ;
    END
  END sram_din_b[22]
  PIN sram_din_b[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 531.120 4.000 531.720 ;
    END
  END sram_din_b[23]
  PIN sram_din_b[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 580.760 1000.000 581.360 ;
    END
  END sram_din_b[24]
  PIN sram_din_b[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 674.450 0.000 674.730 4.000 ;
    END
  END sram_din_b[25]
  PIN sram_din_b[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 673.530 1496.000 673.810 1500.000 ;
    END
  END sram_din_b[26]
  PIN sram_din_b[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 680.890 1496.000 681.170 1500.000 ;
    END
  END sram_din_b[27]
  PIN sram_din_b[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 631.080 4.000 631.680 ;
    END
  END sram_din_b[28]
  PIN sram_din_b[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 719.480 1000.000 720.080 ;
    END
  END sram_din_b[29]
  PIN sram_din_b[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 104.080 1000.000 104.680 ;
    END
  END sram_din_b[2]
  PIN sram_din_b[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 707.570 1496.000 707.850 1500.000 ;
    END
  END sram_din_b[30]
  PIN sram_din_b[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 705.880 4.000 706.480 ;
    END
  END sram_din_b[31]
  PIN sram_din_b[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 459.170 0.000 459.450 4.000 ;
    END
  END sram_din_b[3]
  PIN sram_din_b[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 173.440 1000.000 174.040 ;
    END
  END sram_din_b[4]
  PIN sram_din_b[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 212.880 1000.000 213.480 ;
    END
  END sram_din_b[5]
  PIN sram_din_b[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 481.250 0.000 481.530 4.000 ;
    END
  END sram_din_b[6]
  PIN sram_din_b[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 280.880 4.000 281.480 ;
    END
  END sram_din_b[7]
  PIN sram_din_b[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 312.160 1000.000 312.760 ;
    END
  END sram_din_b[8]
  PIN sram_din_b[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 342.080 1000.000 342.680 ;
    END
  END sram_din_b[9]
  PIN sram_dout_a[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 418.230 0.000 418.510 4.000 ;
    END
  END sram_dout_a[0]
  PIN sram_dout_a[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 518.510 1496.000 518.790 1500.000 ;
    END
  END sram_dout_a[10]
  PIN sram_dout_a[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 537.370 1496.000 537.650 1500.000 ;
    END
  END sram_dout_a[11]
  PIN sram_dout_a[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 545.190 1496.000 545.470 1500.000 ;
    END
  END sram_dout_a[12]
  PIN sram_dout_a[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 372.000 1000.000 372.600 ;
    END
  END sram_dout_a[13]
  PIN sram_dout_a[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 581.530 0.000 581.810 4.000 ;
    END
  END sram_dout_a[14]
  PIN sram_dout_a[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 411.440 1000.000 412.040 ;
    END
  END sram_dout_a[15]
  PIN sram_dout_a[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 593.950 1496.000 594.230 1500.000 ;
    END
  END sram_dout_a[16]
  PIN sram_dout_a[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 461.760 1000.000 462.360 ;
    END
  END sram_dout_a[17]
  PIN sram_dout_a[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 443.400 4.000 444.000 ;
    END
  END sram_dout_a[18]
  PIN sram_dout_a[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 616.950 1496.000 617.230 1500.000 ;
    END
  END sram_dout_a[19]
  PIN sram_dout_a[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 432.950 0.000 433.230 4.000 ;
    END
  END sram_dout_a[1]
  PIN sram_dout_a[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 633.510 0.000 633.790 4.000 ;
    END
  END sram_dout_a[20]
  PIN sram_dout_a[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 632.130 1496.000 632.410 1500.000 ;
    END
  END sram_dout_a[21]
  PIN sram_dout_a[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 643.170 1496.000 643.450 1500.000 ;
    END
  END sram_dout_a[22]
  PIN sram_dout_a[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 663.410 0.000 663.690 4.000 ;
    END
  END sram_dout_a[23]
  PIN sram_dout_a[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 658.350 1496.000 658.630 1500.000 ;
    END
  END sram_dout_a[24]
  PIN sram_dout_a[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 555.600 4.000 556.200 ;
    END
  END sram_dout_a[25]
  PIN sram_dout_a[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 681.810 0.000 682.090 4.000 ;
    END
  END sram_dout_a[26]
  PIN sram_dout_a[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 693.310 0.000 693.590 4.000 ;
    END
  END sram_dout_a[27]
  PIN sram_dout_a[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 692.390 1496.000 692.670 1500.000 ;
    END
  END sram_dout_a[28]
  PIN sram_dout_a[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 696.990 0.000 697.270 4.000 ;
    END
  END sram_dout_a[29]
  PIN sram_dout_a[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 443.990 0.000 444.270 4.000 ;
    END
  END sram_dout_a[2]
  PIN sram_dout_a[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 700.670 0.000 700.950 4.000 ;
    END
  END sram_dout_a[30]
  PIN sram_dout_a[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 708.030 0.000 708.310 4.000 ;
    END
  END sram_dout_a[31]
  PIN sram_dout_a[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 469.750 1496.000 470.030 1500.000 ;
    END
  END sram_dout_a[3]
  PIN sram_dout_a[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 168.000 4.000 168.600 ;
    END
  END sram_dout_a[4]
  PIN sram_dout_a[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 484.930 1496.000 485.210 1500.000 ;
    END
  END sram_dout_a[5]
  PIN sram_dout_a[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 484.930 0.000 485.210 4.000 ;
    END
  END sram_dout_a[6]
  PIN sram_dout_a[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 503.790 0.000 504.070 4.000 ;
    END
  END sram_dout_a[7]
  PIN sram_dout_a[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 322.360 1000.000 322.960 ;
    END
  END sram_dout_a[8]
  PIN sram_dout_a[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 352.280 1000.000 352.880 ;
    END
  END sram_dout_a[9]
  PIN sram_mask_b[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 447.210 1496.000 447.490 1500.000 ;
    END
  END sram_mask_b[0]
  PIN sram_mask_b[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 54.440 1000.000 55.040 ;
    END
  END sram_mask_b[1]
  PIN sram_mask_b[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 113.600 1000.000 114.200 ;
    END
  END sram_mask_b[2]
  PIN sram_mask_b[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 118.360 4.000 118.960 ;
    END
  END sram_mask_b[3]
  PIN sram_web_b
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 432.030 1496.000 432.310 1500.000 ;
    END
  END sram_web_b
  PIN trng_buffer_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 24.520 1000.000 25.120 ;
    END
  END trng_buffer_i[0]
  PIN trng_buffer_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 544.270 0.000 544.550 4.000 ;
    END
  END trng_buffer_i[10]
  PIN trng_buffer_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 361.800 1000.000 362.400 ;
    END
  END trng_buffer_i[11]
  PIN trng_buffer_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 548.870 1496.000 549.150 1500.000 ;
    END
  END trng_buffer_i[12]
  PIN trng_buffer_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 567.730 1496.000 568.010 1500.000 ;
    END
  END trng_buffer_i[13]
  PIN trng_buffer_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 391.720 1000.000 392.320 ;
    END
  END trng_buffer_i[14]
  PIN trng_buffer_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 593.030 0.000 593.310 4.000 ;
    END
  END trng_buffer_i[15]
  PIN trng_buffer_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 598.090 1496.000 598.370 1500.000 ;
    END
  END trng_buffer_i[16]
  PIN trng_buffer_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 601.770 1496.000 602.050 1500.000 ;
    END
  END trng_buffer_i[17]
  PIN trng_buffer_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 455.640 4.000 456.240 ;
    END
  END trng_buffer_i[18]
  PIN trng_buffer_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 468.560 4.000 469.160 ;
    END
  END trng_buffer_i[19]
  PIN trng_buffer_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 63.960 1000.000 64.560 ;
    END
  END trng_buffer_i[1]
  PIN trng_buffer_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 480.800 4.000 481.400 ;
    END
  END trng_buffer_i[20]
  PIN trng_buffer_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 505.960 4.000 506.560 ;
    END
  END trng_buffer_i[21]
  PIN trng_buffer_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 646.850 1496.000 647.130 1500.000 ;
    END
  END trng_buffer_i[22]
  PIN trng_buffer_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 550.840 1000.000 551.440 ;
    END
  END trng_buffer_i[23]
  PIN trng_buffer_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 590.280 1000.000 590.880 ;
    END
  END trng_buffer_i[24]
  PIN trng_buffer_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 678.130 0.000 678.410 4.000 ;
    END
  END trng_buffer_i[25]
  PIN trng_buffer_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 685.950 0.000 686.230 4.000 ;
    END
  END trng_buffer_i[26]
  PIN trng_buffer_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 684.570 1496.000 684.850 1500.000 ;
    END
  END trng_buffer_i[27]
  PIN trng_buffer_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 643.320 4.000 643.920 ;
    END
  END trng_buffer_i[28]
  PIN trng_buffer_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 668.480 4.000 669.080 ;
    END
  END trng_buffer_i[29]
  PIN trng_buffer_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 461.930 1496.000 462.210 1500.000 ;
    END
  END trng_buffer_i[2]
  PIN trng_buffer_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 704.350 0.000 704.630 4.000 ;
    END
  END trng_buffer_i[30]
  PIN trng_buffer_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 759.600 1000.000 760.200 ;
    END
  END trng_buffer_i[31]
  PIN trng_buffer_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 153.720 1000.000 154.320 ;
    END
  END trng_buffer_i[3]
  PIN trng_buffer_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 470.210 0.000 470.490 4.000 ;
    END
  END trng_buffer_i[4]
  PIN trng_buffer_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 223.080 1000.000 223.680 ;
    END
  END trng_buffer_i[5]
  PIN trng_buffer_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 488.610 0.000 488.890 4.000 ;
    END
  END trng_buffer_i[6]
  PIN trng_buffer_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 507.470 0.000 507.750 4.000 ;
    END
  END trng_buffer_i[7]
  PIN trng_buffer_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 332.560 1000.000 333.160 ;
    END
  END trng_buffer_i[8]
  PIN trng_buffer_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 503.790 1496.000 504.070 1500.000 ;
    END
  END trng_buffer_i[9]
  PIN trng_wb_ack_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 410.410 0.000 410.690 4.000 ;
    END
  END trng_wb_ack_i
  PIN trng_wb_adr_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 55.800 4.000 56.400 ;
    END
  END trng_wb_adr_o[0]
  PIN trng_wb_adr_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 454.570 1496.000 454.850 1500.000 ;
    END
  END trng_wb_adr_o[1]
  PIN trng_wb_adr_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 123.800 1000.000 124.400 ;
    END
  END trng_wb_adr_o[2]
  PIN trng_wb_adr_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 462.850 0.000 463.130 4.000 ;
    END
  END trng_wb_adr_o[3]
  PIN trng_wb_adr_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 182.960 1000.000 183.560 ;
    END
  END trng_wb_adr_o[4]
  PIN trng_wb_adr_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 218.320 4.000 218.920 ;
    END
  END trng_wb_adr_o[5]
  PIN trng_wb_adr_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 255.720 4.000 256.320 ;
    END
  END trng_wb_adr_o[6]
  PIN trng_wb_adr_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 293.120 4.000 293.720 ;
    END
  END trng_wb_adr_o[7]
  PIN trng_wb_adr_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 518.510 0.000 518.790 4.000 ;
    END
  END trng_wb_adr_o[8]
  PIN trng_wb_cyc_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 435.710 1496.000 435.990 1500.000 ;
    END
  END trng_wb_cyc_o
  PIN trng_wb_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.040 4.000 68.640 ;
    END
  END trng_wb_dat_i[0]
  PIN trng_wb_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 522.650 1496.000 522.930 1500.000 ;
    END
  END trng_wb_dat_i[10]
  PIN trng_wb_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 552.090 0.000 552.370 4.000 ;
    END
  END trng_wb_dat_i[11]
  PIN trng_wb_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 552.550 1496.000 552.830 1500.000 ;
    END
  END trng_wb_dat_i[12]
  PIN trng_wb_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 574.170 0.000 574.450 4.000 ;
    END
  END trng_wb_dat_i[13]
  PIN trng_wb_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 579.230 1496.000 579.510 1500.000 ;
    END
  END trng_wb_dat_i[14]
  PIN trng_wb_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 586.590 1496.000 586.870 1500.000 ;
    END
  END trng_wb_dat_i[15]
  PIN trng_wb_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 406.000 4.000 406.600 ;
    END
  END trng_wb_dat_i[16]
  PIN trng_wb_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 605.450 1496.000 605.730 1500.000 ;
    END
  END trng_wb_dat_i[17]
  PIN trng_wb_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 613.270 1496.000 613.550 1500.000 ;
    END
  END trng_wb_dat_i[18]
  PIN trng_wb_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 491.000 1000.000 491.600 ;
    END
  END trng_wb_dat_i[19]
  PIN trng_wb_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 74.160 1000.000 74.760 ;
    END
  END trng_wb_dat_i[1]
  PIN trng_wb_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 637.190 0.000 637.470 4.000 ;
    END
  END trng_wb_dat_i[20]
  PIN trng_wb_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 635.810 1496.000 636.090 1500.000 ;
    END
  END trng_wb_dat_i[21]
  PIN trng_wb_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 540.640 1000.000 541.240 ;
    END
  END trng_wb_dat_i[22]
  PIN trng_wb_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 561.040 1000.000 561.640 ;
    END
  END trng_wb_dat_i[23]
  PIN trng_wb_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 662.030 1496.000 662.310 1500.000 ;
    END
  END trng_wb_dat_i[24]
  PIN trng_wb_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 665.710 1496.000 665.990 1500.000 ;
    END
  END trng_wb_dat_i[25]
  PIN trng_wb_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 689.630 0.000 689.910 4.000 ;
    END
  END trng_wb_dat_i[26]
  PIN trng_wb_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 660.320 1000.000 660.920 ;
    END
  END trng_wb_dat_i[27]
  PIN trng_wb_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 680.040 1000.000 680.640 ;
    END
  END trng_wb_dat_i[28]
  PIN trng_wb_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 696.070 1496.000 696.350 1500.000 ;
    END
  END trng_wb_dat_i[29]
  PIN trng_wb_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 106.120 4.000 106.720 ;
    END
  END trng_wb_dat_i[2]
  PIN trng_wb_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 739.880 1000.000 740.480 ;
    END
  END trng_wb_dat_i[30]
  PIN trng_wb_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 711.710 0.000 711.990 4.000 ;
    END
  END trng_wb_dat_i[31]
  PIN trng_wb_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 163.240 1000.000 163.840 ;
    END
  END trng_wb_dat_i[3]
  PIN trng_wb_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 180.920 4.000 181.520 ;
    END
  END trng_wb_dat_i[4]
  PIN trng_wb_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 477.570 0.000 477.850 4.000 ;
    END
  END trng_wb_dat_i[5]
  PIN trng_wb_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 492.290 0.000 492.570 4.000 ;
    END
  END trng_wb_dat_i[6]
  PIN trng_wb_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 282.920 1000.000 283.520 ;
    END
  END trng_wb_dat_i[7]
  PIN trng_wb_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 522.190 0.000 522.470 4.000 ;
    END
  END trng_wb_dat_i[8]
  PIN trng_wb_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 507.470 1496.000 507.750 1500.000 ;
    END
  END trng_wb_dat_i[9]
  PIN trng_wb_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 450.890 1496.000 451.170 1500.000 ;
    END
  END trng_wb_dat_o[0]
  PIN trng_wb_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 548.410 0.000 548.690 4.000 ;
    END
  END trng_wb_dat_o[10]
  PIN trng_wb_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 555.770 0.000 556.050 4.000 ;
    END
  END trng_wb_dat_o[11]
  PIN trng_wb_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 566.810 0.000 567.090 4.000 ;
    END
  END trng_wb_dat_o[12]
  PIN trng_wb_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 382.200 1000.000 382.800 ;
    END
  END trng_wb_dat_o[13]
  PIN trng_wb_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 585.210 0.000 585.490 4.000 ;
    END
  END trng_wb_dat_o[14]
  PIN trng_wb_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 596.710 0.000 596.990 4.000 ;
    END
  END trng_wb_dat_o[15]
  PIN trng_wb_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 421.640 1000.000 422.240 ;
    END
  END trng_wb_dat_o[16]
  PIN trng_wb_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 471.280 1000.000 471.880 ;
    END
  END trng_wb_dat_o[17]
  PIN trng_wb_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 611.430 0.000 611.710 4.000 ;
    END
  END trng_wb_dat_o[18]
  PIN trng_wb_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 620.630 1496.000 620.910 1500.000 ;
    END
  END trng_wb_dat_o[19]
  PIN trng_wb_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 83.680 1000.000 84.280 ;
    END
  END trng_wb_dat_o[1]
  PIN trng_wb_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 641.330 0.000 641.610 4.000 ;
    END
  END trng_wb_dat_o[20]
  PIN trng_wb_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 648.690 0.000 648.970 4.000 ;
    END
  END trng_wb_dat_o[21]
  PIN trng_wb_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 650.990 1496.000 651.270 1500.000 ;
    END
  END trng_wb_dat_o[22]
  PIN trng_wb_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 667.090 0.000 667.370 4.000 ;
    END
  END trng_wb_dat_o[23]
  PIN trng_wb_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 600.480 1000.000 601.080 ;
    END
  END trng_wb_dat_o[24]
  PIN trng_wb_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 568.520 4.000 569.120 ;
    END
  END trng_wb_dat_o[25]
  PIN trng_wb_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 677.210 1496.000 677.490 1500.000 ;
    END
  END trng_wb_dat_o[26]
  PIN trng_wb_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 669.840 1000.000 670.440 ;
    END
  END trng_wb_dat_o[27]
  PIN trng_wb_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 655.560 4.000 656.160 ;
    END
  END trng_wb_dat_o[28]
  PIN trng_wb_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 680.720 4.000 681.320 ;
    END
  END trng_wb_dat_o[29]
  PIN trng_wb_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 447.670 0.000 447.950 4.000 ;
    END
  END trng_wb_dat_o[2]
  PIN trng_wb_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 693.640 4.000 694.240 ;
    END
  END trng_wb_dat_o[30]
  PIN trng_wb_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 715.390 0.000 715.670 4.000 ;
    END
  END trng_wb_dat_o[31]
  PIN trng_wb_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 473.430 1496.000 473.710 1500.000 ;
    END
  END trng_wb_dat_o[3]
  PIN trng_wb_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 193.160 4.000 193.760 ;
    END
  END trng_wb_dat_o[4]
  PIN trng_wb_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 233.280 1000.000 233.880 ;
    END
  END trng_wb_dat_o[5]
  PIN trng_wb_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 488.610 1496.000 488.890 1500.000 ;
    END
  END trng_wb_dat_o[6]
  PIN trng_wb_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 292.440 1000.000 293.040 ;
    END
  END trng_wb_dat_o[7]
  PIN trng_wb_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 525.870 0.000 526.150 4.000 ;
    END
  END trng_wb_dat_o[8]
  PIN trng_wb_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 511.150 1496.000 511.430 1500.000 ;
    END
  END trng_wb_dat_o[9]
  PIN trng_wb_stb_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 439.390 1496.000 439.670 1500.000 ;
    END
  END trng_wb_stb_o
  PIN trng_wb_we_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 443.070 1496.000 443.350 1500.000 ;
    END
  END trng_wb_we_o
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 942.640 10.640 944.240 1488.080 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 865.840 10.640 867.440 1488.080 ;
    END
  END vssd1
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.930 0.000 2.210 4.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.610 0.000 5.890 4.000 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.290 0.000 9.570 4.000 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.010 0.000 24.290 4.000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.510 0.000 150.790 4.000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.550 0.000 161.830 4.000 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 172.590 0.000 172.870 4.000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 184.090 0.000 184.370 4.000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 195.130 0.000 195.410 4.000 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 206.170 0.000 206.450 4.000 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 217.210 0.000 217.490 4.000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 228.250 0.000 228.530 4.000 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 239.750 0.000 240.030 4.000 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 250.790 0.000 251.070 4.000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.730 0.000 39.010 4.000 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 261.830 0.000 262.110 4.000 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 272.870 0.000 273.150 4.000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 284.370 0.000 284.650 4.000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 295.410 0.000 295.690 4.000 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 306.450 0.000 306.730 4.000 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 317.490 0.000 317.770 4.000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 328.990 0.000 329.270 4.000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 340.030 0.000 340.310 4.000 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 351.070 0.000 351.350 4.000 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 362.110 0.000 362.390 4.000 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.910 0.000 54.190 4.000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 373.610 0.000 373.890 4.000 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 384.650 0.000 384.930 4.000 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.630 0.000 68.910 4.000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.350 0.000 83.630 4.000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.850 0.000 95.130 4.000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 105.890 0.000 106.170 4.000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.930 0.000 117.210 4.000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.970 0.000 128.250 4.000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.470 0.000 139.750 4.000 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.970 0.000 13.250 4.000 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.690 0.000 27.970 4.000 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 154.190 0.000 154.470 4.000 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 165.230 0.000 165.510 4.000 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 176.270 0.000 176.550 4.000 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 187.770 0.000 188.050 4.000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 198.810 0.000 199.090 4.000 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.850 0.000 210.130 4.000 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 220.890 0.000 221.170 4.000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 232.390 0.000 232.670 4.000 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 243.430 0.000 243.710 4.000 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.470 0.000 254.750 4.000 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.410 0.000 42.690 4.000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 265.510 0.000 265.790 4.000 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 277.010 0.000 277.290 4.000 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 288.050 0.000 288.330 4.000 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 299.090 0.000 299.370 4.000 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 310.130 0.000 310.410 4.000 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 321.630 0.000 321.910 4.000 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 332.670 0.000 332.950 4.000 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 343.710 0.000 343.990 4.000 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 354.750 0.000 355.030 4.000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 366.250 0.000 366.530 4.000 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.590 0.000 57.870 4.000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 377.290 0.000 377.570 4.000 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 388.330 0.000 388.610 4.000 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.310 0.000 72.590 4.000 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.030 0.000 87.310 4.000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.530 0.000 98.810 4.000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.570 0.000 109.850 4.000 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.610 0.000 120.890 4.000 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 131.650 0.000 131.930 4.000 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 143.150 0.000 143.430 4.000 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.370 0.000 31.650 4.000 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.870 0.000 158.150 4.000 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 168.910 0.000 169.190 4.000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.950 0.000 180.230 4.000 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 191.450 0.000 191.730 4.000 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.490 0.000 202.770 4.000 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 213.530 0.000 213.810 4.000 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 224.570 0.000 224.850 4.000 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 236.070 0.000 236.350 4.000 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 247.110 0.000 247.390 4.000 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 258.150 0.000 258.430 4.000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.090 0.000 46.370 4.000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 269.190 0.000 269.470 4.000 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 280.690 0.000 280.970 4.000 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 291.730 0.000 292.010 4.000 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 302.770 0.000 303.050 4.000 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 313.810 0.000 314.090 4.000 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 325.310 0.000 325.590 4.000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 336.350 0.000 336.630 4.000 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 347.390 0.000 347.670 4.000 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 358.430 0.000 358.710 4.000 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 369.930 0.000 370.210 4.000 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.270 0.000 61.550 4.000 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 380.970 0.000 381.250 4.000 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 392.010 0.000 392.290 4.000 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.990 0.000 76.270 4.000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.710 0.000 90.990 4.000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.210 0.000 102.490 4.000 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 113.250 0.000 113.530 4.000 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 124.290 0.000 124.570 4.000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.330 0.000 135.610 4.000 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 146.830 0.000 147.110 4.000 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.050 0.000 35.330 4.000 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.230 0.000 50.510 4.000 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.950 0.000 65.230 4.000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.670 0.000 79.950 4.000 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.650 0.000 16.930 4.000 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.330 0.000 20.610 4.000 ;
    END
  END wbs_we_i
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 994.060 1487.925 ;
      LAYER met1 ;
        RECT 1.910 4.460 997.670 1488.080 ;
      LAYER met2 ;
        RECT 2.490 1495.720 5.330 1496.410 ;
        RECT 6.170 1495.720 9.010 1496.410 ;
        RECT 9.850 1495.720 12.690 1496.410 ;
        RECT 13.530 1495.720 16.370 1496.410 ;
        RECT 17.210 1495.720 20.510 1496.410 ;
        RECT 21.350 1495.720 24.190 1496.410 ;
        RECT 25.030 1495.720 27.870 1496.410 ;
        RECT 28.710 1495.720 31.550 1496.410 ;
        RECT 32.390 1495.720 35.230 1496.410 ;
        RECT 36.070 1495.720 39.370 1496.410 ;
        RECT 40.210 1495.720 43.050 1496.410 ;
        RECT 43.890 1495.720 46.730 1496.410 ;
        RECT 47.570 1495.720 50.410 1496.410 ;
        RECT 51.250 1495.720 54.090 1496.410 ;
        RECT 54.930 1495.720 58.230 1496.410 ;
        RECT 59.070 1495.720 61.910 1496.410 ;
        RECT 62.750 1495.720 65.590 1496.410 ;
        RECT 66.430 1495.720 69.270 1496.410 ;
        RECT 70.110 1495.720 72.950 1496.410 ;
        RECT 73.790 1495.720 77.090 1496.410 ;
        RECT 77.930 1495.720 80.770 1496.410 ;
        RECT 81.610 1495.720 84.450 1496.410 ;
        RECT 85.290 1495.720 88.130 1496.410 ;
        RECT 88.970 1495.720 91.810 1496.410 ;
        RECT 92.650 1495.720 95.950 1496.410 ;
        RECT 96.790 1495.720 99.630 1496.410 ;
        RECT 100.470 1495.720 103.310 1496.410 ;
        RECT 104.150 1495.720 106.990 1496.410 ;
        RECT 107.830 1495.720 110.670 1496.410 ;
        RECT 111.510 1495.720 114.810 1496.410 ;
        RECT 115.650 1495.720 118.490 1496.410 ;
        RECT 119.330 1495.720 122.170 1496.410 ;
        RECT 123.010 1495.720 125.850 1496.410 ;
        RECT 126.690 1495.720 129.530 1496.410 ;
        RECT 130.370 1495.720 133.670 1496.410 ;
        RECT 134.510 1495.720 137.350 1496.410 ;
        RECT 138.190 1495.720 141.030 1496.410 ;
        RECT 141.870 1495.720 144.710 1496.410 ;
        RECT 145.550 1495.720 148.390 1496.410 ;
        RECT 149.230 1495.720 152.530 1496.410 ;
        RECT 153.370 1495.720 156.210 1496.410 ;
        RECT 157.050 1495.720 159.890 1496.410 ;
        RECT 160.730 1495.720 163.570 1496.410 ;
        RECT 164.410 1495.720 167.250 1496.410 ;
        RECT 168.090 1495.720 171.390 1496.410 ;
        RECT 172.230 1495.720 175.070 1496.410 ;
        RECT 175.910 1495.720 178.750 1496.410 ;
        RECT 179.590 1495.720 182.430 1496.410 ;
        RECT 183.270 1495.720 186.110 1496.410 ;
        RECT 186.950 1495.720 190.250 1496.410 ;
        RECT 191.090 1495.720 193.930 1496.410 ;
        RECT 194.770 1495.720 197.610 1496.410 ;
        RECT 198.450 1495.720 201.290 1496.410 ;
        RECT 202.130 1495.720 205.430 1496.410 ;
        RECT 206.270 1495.720 209.110 1496.410 ;
        RECT 209.950 1495.720 212.790 1496.410 ;
        RECT 213.630 1495.720 216.470 1496.410 ;
        RECT 217.310 1495.720 220.150 1496.410 ;
        RECT 220.990 1495.720 224.290 1496.410 ;
        RECT 225.130 1495.720 227.970 1496.410 ;
        RECT 228.810 1495.720 231.650 1496.410 ;
        RECT 232.490 1495.720 235.330 1496.410 ;
        RECT 236.170 1495.720 239.010 1496.410 ;
        RECT 239.850 1495.720 243.150 1496.410 ;
        RECT 243.990 1495.720 246.830 1496.410 ;
        RECT 247.670 1495.720 250.510 1496.410 ;
        RECT 251.350 1495.720 254.190 1496.410 ;
        RECT 255.030 1495.720 257.870 1496.410 ;
        RECT 258.710 1495.720 262.010 1496.410 ;
        RECT 262.850 1495.720 265.690 1496.410 ;
        RECT 266.530 1495.720 269.370 1496.410 ;
        RECT 270.210 1495.720 273.050 1496.410 ;
        RECT 273.890 1495.720 276.730 1496.410 ;
        RECT 277.570 1495.720 280.870 1496.410 ;
        RECT 281.710 1495.720 284.550 1496.410 ;
        RECT 285.390 1495.720 288.230 1496.410 ;
        RECT 289.070 1495.720 291.910 1496.410 ;
        RECT 292.750 1495.720 295.590 1496.410 ;
        RECT 296.430 1495.720 299.730 1496.410 ;
        RECT 300.570 1495.720 303.410 1496.410 ;
        RECT 304.250 1495.720 307.090 1496.410 ;
        RECT 307.930 1495.720 310.770 1496.410 ;
        RECT 311.610 1495.720 314.450 1496.410 ;
        RECT 315.290 1495.720 318.590 1496.410 ;
        RECT 319.430 1495.720 322.270 1496.410 ;
        RECT 323.110 1495.720 325.950 1496.410 ;
        RECT 326.790 1495.720 329.630 1496.410 ;
        RECT 330.470 1495.720 333.310 1496.410 ;
        RECT 334.150 1495.720 337.450 1496.410 ;
        RECT 338.290 1495.720 341.130 1496.410 ;
        RECT 341.970 1495.720 344.810 1496.410 ;
        RECT 345.650 1495.720 348.490 1496.410 ;
        RECT 349.330 1495.720 352.170 1496.410 ;
        RECT 353.010 1495.720 356.310 1496.410 ;
        RECT 357.150 1495.720 359.990 1496.410 ;
        RECT 360.830 1495.720 363.670 1496.410 ;
        RECT 364.510 1495.720 367.350 1496.410 ;
        RECT 368.190 1495.720 371.030 1496.410 ;
        RECT 371.870 1495.720 375.170 1496.410 ;
        RECT 376.010 1495.720 378.850 1496.410 ;
        RECT 379.690 1495.720 382.530 1496.410 ;
        RECT 383.370 1495.720 386.210 1496.410 ;
        RECT 387.050 1495.720 389.890 1496.410 ;
        RECT 390.730 1495.720 394.030 1496.410 ;
        RECT 394.870 1495.720 397.710 1496.410 ;
        RECT 398.550 1495.720 401.390 1496.410 ;
        RECT 402.230 1495.720 405.070 1496.410 ;
        RECT 405.910 1495.720 409.210 1496.410 ;
        RECT 410.050 1495.720 412.890 1496.410 ;
        RECT 413.730 1495.720 416.570 1496.410 ;
        RECT 417.410 1495.720 420.250 1496.410 ;
        RECT 421.090 1495.720 423.930 1496.410 ;
        RECT 424.770 1495.720 428.070 1496.410 ;
        RECT 428.910 1495.720 431.750 1496.410 ;
        RECT 432.590 1495.720 435.430 1496.410 ;
        RECT 436.270 1495.720 439.110 1496.410 ;
        RECT 439.950 1495.720 442.790 1496.410 ;
        RECT 443.630 1495.720 446.930 1496.410 ;
        RECT 447.770 1495.720 450.610 1496.410 ;
        RECT 451.450 1495.720 454.290 1496.410 ;
        RECT 455.130 1495.720 457.970 1496.410 ;
        RECT 458.810 1495.720 461.650 1496.410 ;
        RECT 462.490 1495.720 465.790 1496.410 ;
        RECT 466.630 1495.720 469.470 1496.410 ;
        RECT 470.310 1495.720 473.150 1496.410 ;
        RECT 473.990 1495.720 476.830 1496.410 ;
        RECT 477.670 1495.720 480.510 1496.410 ;
        RECT 481.350 1495.720 484.650 1496.410 ;
        RECT 485.490 1495.720 488.330 1496.410 ;
        RECT 489.170 1495.720 492.010 1496.410 ;
        RECT 492.850 1495.720 495.690 1496.410 ;
        RECT 496.530 1495.720 499.370 1496.410 ;
        RECT 500.210 1495.720 503.510 1496.410 ;
        RECT 504.350 1495.720 507.190 1496.410 ;
        RECT 508.030 1495.720 510.870 1496.410 ;
        RECT 511.710 1495.720 514.550 1496.410 ;
        RECT 515.390 1495.720 518.230 1496.410 ;
        RECT 519.070 1495.720 522.370 1496.410 ;
        RECT 523.210 1495.720 526.050 1496.410 ;
        RECT 526.890 1495.720 529.730 1496.410 ;
        RECT 530.570 1495.720 533.410 1496.410 ;
        RECT 534.250 1495.720 537.090 1496.410 ;
        RECT 537.930 1495.720 541.230 1496.410 ;
        RECT 542.070 1495.720 544.910 1496.410 ;
        RECT 545.750 1495.720 548.590 1496.410 ;
        RECT 549.430 1495.720 552.270 1496.410 ;
        RECT 553.110 1495.720 555.950 1496.410 ;
        RECT 556.790 1495.720 560.090 1496.410 ;
        RECT 560.930 1495.720 563.770 1496.410 ;
        RECT 564.610 1495.720 567.450 1496.410 ;
        RECT 568.290 1495.720 571.130 1496.410 ;
        RECT 571.970 1495.720 574.810 1496.410 ;
        RECT 575.650 1495.720 578.950 1496.410 ;
        RECT 579.790 1495.720 582.630 1496.410 ;
        RECT 583.470 1495.720 586.310 1496.410 ;
        RECT 587.150 1495.720 589.990 1496.410 ;
        RECT 590.830 1495.720 593.670 1496.410 ;
        RECT 594.510 1495.720 597.810 1496.410 ;
        RECT 598.650 1495.720 601.490 1496.410 ;
        RECT 602.330 1495.720 605.170 1496.410 ;
        RECT 606.010 1495.720 608.850 1496.410 ;
        RECT 609.690 1495.720 612.990 1496.410 ;
        RECT 613.830 1495.720 616.670 1496.410 ;
        RECT 617.510 1495.720 620.350 1496.410 ;
        RECT 621.190 1495.720 624.030 1496.410 ;
        RECT 624.870 1495.720 627.710 1496.410 ;
        RECT 628.550 1495.720 631.850 1496.410 ;
        RECT 632.690 1495.720 635.530 1496.410 ;
        RECT 636.370 1495.720 639.210 1496.410 ;
        RECT 640.050 1495.720 642.890 1496.410 ;
        RECT 643.730 1495.720 646.570 1496.410 ;
        RECT 647.410 1495.720 650.710 1496.410 ;
        RECT 651.550 1495.720 654.390 1496.410 ;
        RECT 655.230 1495.720 658.070 1496.410 ;
        RECT 658.910 1495.720 661.750 1496.410 ;
        RECT 662.590 1495.720 665.430 1496.410 ;
        RECT 666.270 1495.720 669.570 1496.410 ;
        RECT 670.410 1495.720 673.250 1496.410 ;
        RECT 674.090 1495.720 676.930 1496.410 ;
        RECT 677.770 1495.720 680.610 1496.410 ;
        RECT 681.450 1495.720 684.290 1496.410 ;
        RECT 685.130 1495.720 688.430 1496.410 ;
        RECT 689.270 1495.720 692.110 1496.410 ;
        RECT 692.950 1495.720 695.790 1496.410 ;
        RECT 696.630 1495.720 699.470 1496.410 ;
        RECT 700.310 1495.720 703.150 1496.410 ;
        RECT 703.990 1495.720 707.290 1496.410 ;
        RECT 708.130 1495.720 710.970 1496.410 ;
        RECT 711.810 1495.720 714.650 1496.410 ;
        RECT 715.490 1495.720 718.330 1496.410 ;
        RECT 719.170 1495.720 722.010 1496.410 ;
        RECT 722.850 1495.720 726.150 1496.410 ;
        RECT 726.990 1495.720 729.830 1496.410 ;
        RECT 730.670 1495.720 733.510 1496.410 ;
        RECT 734.350 1495.720 737.190 1496.410 ;
        RECT 738.030 1495.720 740.870 1496.410 ;
        RECT 741.710 1495.720 745.010 1496.410 ;
        RECT 745.850 1495.720 748.690 1496.410 ;
        RECT 749.530 1495.720 752.370 1496.410 ;
        RECT 753.210 1495.720 756.050 1496.410 ;
        RECT 756.890 1495.720 759.730 1496.410 ;
        RECT 760.570 1495.720 763.870 1496.410 ;
        RECT 764.710 1495.720 767.550 1496.410 ;
        RECT 768.390 1495.720 771.230 1496.410 ;
        RECT 772.070 1495.720 774.910 1496.410 ;
        RECT 775.750 1495.720 778.590 1496.410 ;
        RECT 779.430 1495.720 782.730 1496.410 ;
        RECT 783.570 1495.720 786.410 1496.410 ;
        RECT 787.250 1495.720 790.090 1496.410 ;
        RECT 790.930 1495.720 793.770 1496.410 ;
        RECT 794.610 1495.720 797.450 1496.410 ;
        RECT 798.290 1495.720 801.590 1496.410 ;
        RECT 802.430 1495.720 805.270 1496.410 ;
        RECT 806.110 1495.720 808.950 1496.410 ;
        RECT 809.790 1495.720 812.630 1496.410 ;
        RECT 813.470 1495.720 816.770 1496.410 ;
        RECT 817.610 1495.720 820.450 1496.410 ;
        RECT 821.290 1495.720 824.130 1496.410 ;
        RECT 824.970 1495.720 827.810 1496.410 ;
        RECT 828.650 1495.720 831.490 1496.410 ;
        RECT 832.330 1495.720 835.630 1496.410 ;
        RECT 836.470 1495.720 839.310 1496.410 ;
        RECT 840.150 1495.720 842.990 1496.410 ;
        RECT 843.830 1495.720 846.670 1496.410 ;
        RECT 847.510 1495.720 850.350 1496.410 ;
        RECT 851.190 1495.720 854.490 1496.410 ;
        RECT 855.330 1495.720 858.170 1496.410 ;
        RECT 859.010 1495.720 861.850 1496.410 ;
        RECT 862.690 1495.720 865.530 1496.410 ;
        RECT 866.370 1495.720 869.210 1496.410 ;
        RECT 870.050 1495.720 873.350 1496.410 ;
        RECT 874.190 1495.720 877.030 1496.410 ;
        RECT 877.870 1495.720 880.710 1496.410 ;
        RECT 881.550 1495.720 884.390 1496.410 ;
        RECT 885.230 1495.720 888.070 1496.410 ;
        RECT 888.910 1495.720 892.210 1496.410 ;
        RECT 893.050 1495.720 895.890 1496.410 ;
        RECT 896.730 1495.720 899.570 1496.410 ;
        RECT 900.410 1495.720 903.250 1496.410 ;
        RECT 904.090 1495.720 906.930 1496.410 ;
        RECT 907.770 1495.720 911.070 1496.410 ;
        RECT 911.910 1495.720 914.750 1496.410 ;
        RECT 915.590 1495.720 918.430 1496.410 ;
        RECT 919.270 1495.720 922.110 1496.410 ;
        RECT 922.950 1495.720 925.790 1496.410 ;
        RECT 926.630 1495.720 929.930 1496.410 ;
        RECT 930.770 1495.720 933.610 1496.410 ;
        RECT 934.450 1495.720 937.290 1496.410 ;
        RECT 938.130 1495.720 940.970 1496.410 ;
        RECT 941.810 1495.720 944.650 1496.410 ;
        RECT 945.490 1495.720 948.790 1496.410 ;
        RECT 949.630 1495.720 952.470 1496.410 ;
        RECT 953.310 1495.720 956.150 1496.410 ;
        RECT 956.990 1495.720 959.830 1496.410 ;
        RECT 960.670 1495.720 963.510 1496.410 ;
        RECT 964.350 1495.720 967.650 1496.410 ;
        RECT 968.490 1495.720 971.330 1496.410 ;
        RECT 972.170 1495.720 975.010 1496.410 ;
        RECT 975.850 1495.720 978.690 1496.410 ;
        RECT 979.530 1495.720 982.370 1496.410 ;
        RECT 983.210 1495.720 986.510 1496.410 ;
        RECT 987.350 1495.720 990.190 1496.410 ;
        RECT 991.030 1495.720 993.870 1496.410 ;
        RECT 994.710 1495.720 997.550 1496.410 ;
        RECT 1.940 4.280 997.640 1495.720 ;
        RECT 2.490 3.670 5.330 4.280 ;
        RECT 6.170 3.670 9.010 4.280 ;
        RECT 9.850 3.670 12.690 4.280 ;
        RECT 13.530 3.670 16.370 4.280 ;
        RECT 17.210 3.670 20.050 4.280 ;
        RECT 20.890 3.670 23.730 4.280 ;
        RECT 24.570 3.670 27.410 4.280 ;
        RECT 28.250 3.670 31.090 4.280 ;
        RECT 31.930 3.670 34.770 4.280 ;
        RECT 35.610 3.670 38.450 4.280 ;
        RECT 39.290 3.670 42.130 4.280 ;
        RECT 42.970 3.670 45.810 4.280 ;
        RECT 46.650 3.670 49.950 4.280 ;
        RECT 50.790 3.670 53.630 4.280 ;
        RECT 54.470 3.670 57.310 4.280 ;
        RECT 58.150 3.670 60.990 4.280 ;
        RECT 61.830 3.670 64.670 4.280 ;
        RECT 65.510 3.670 68.350 4.280 ;
        RECT 69.190 3.670 72.030 4.280 ;
        RECT 72.870 3.670 75.710 4.280 ;
        RECT 76.550 3.670 79.390 4.280 ;
        RECT 80.230 3.670 83.070 4.280 ;
        RECT 83.910 3.670 86.750 4.280 ;
        RECT 87.590 3.670 90.430 4.280 ;
        RECT 91.270 3.670 94.570 4.280 ;
        RECT 95.410 3.670 98.250 4.280 ;
        RECT 99.090 3.670 101.930 4.280 ;
        RECT 102.770 3.670 105.610 4.280 ;
        RECT 106.450 3.670 109.290 4.280 ;
        RECT 110.130 3.670 112.970 4.280 ;
        RECT 113.810 3.670 116.650 4.280 ;
        RECT 117.490 3.670 120.330 4.280 ;
        RECT 121.170 3.670 124.010 4.280 ;
        RECT 124.850 3.670 127.690 4.280 ;
        RECT 128.530 3.670 131.370 4.280 ;
        RECT 132.210 3.670 135.050 4.280 ;
        RECT 135.890 3.670 139.190 4.280 ;
        RECT 140.030 3.670 142.870 4.280 ;
        RECT 143.710 3.670 146.550 4.280 ;
        RECT 147.390 3.670 150.230 4.280 ;
        RECT 151.070 3.670 153.910 4.280 ;
        RECT 154.750 3.670 157.590 4.280 ;
        RECT 158.430 3.670 161.270 4.280 ;
        RECT 162.110 3.670 164.950 4.280 ;
        RECT 165.790 3.670 168.630 4.280 ;
        RECT 169.470 3.670 172.310 4.280 ;
        RECT 173.150 3.670 175.990 4.280 ;
        RECT 176.830 3.670 179.670 4.280 ;
        RECT 180.510 3.670 183.810 4.280 ;
        RECT 184.650 3.670 187.490 4.280 ;
        RECT 188.330 3.670 191.170 4.280 ;
        RECT 192.010 3.670 194.850 4.280 ;
        RECT 195.690 3.670 198.530 4.280 ;
        RECT 199.370 3.670 202.210 4.280 ;
        RECT 203.050 3.670 205.890 4.280 ;
        RECT 206.730 3.670 209.570 4.280 ;
        RECT 210.410 3.670 213.250 4.280 ;
        RECT 214.090 3.670 216.930 4.280 ;
        RECT 217.770 3.670 220.610 4.280 ;
        RECT 221.450 3.670 224.290 4.280 ;
        RECT 225.130 3.670 227.970 4.280 ;
        RECT 228.810 3.670 232.110 4.280 ;
        RECT 232.950 3.670 235.790 4.280 ;
        RECT 236.630 3.670 239.470 4.280 ;
        RECT 240.310 3.670 243.150 4.280 ;
        RECT 243.990 3.670 246.830 4.280 ;
        RECT 247.670 3.670 250.510 4.280 ;
        RECT 251.350 3.670 254.190 4.280 ;
        RECT 255.030 3.670 257.870 4.280 ;
        RECT 258.710 3.670 261.550 4.280 ;
        RECT 262.390 3.670 265.230 4.280 ;
        RECT 266.070 3.670 268.910 4.280 ;
        RECT 269.750 3.670 272.590 4.280 ;
        RECT 273.430 3.670 276.730 4.280 ;
        RECT 277.570 3.670 280.410 4.280 ;
        RECT 281.250 3.670 284.090 4.280 ;
        RECT 284.930 3.670 287.770 4.280 ;
        RECT 288.610 3.670 291.450 4.280 ;
        RECT 292.290 3.670 295.130 4.280 ;
        RECT 295.970 3.670 298.810 4.280 ;
        RECT 299.650 3.670 302.490 4.280 ;
        RECT 303.330 3.670 306.170 4.280 ;
        RECT 307.010 3.670 309.850 4.280 ;
        RECT 310.690 3.670 313.530 4.280 ;
        RECT 314.370 3.670 317.210 4.280 ;
        RECT 318.050 3.670 321.350 4.280 ;
        RECT 322.190 3.670 325.030 4.280 ;
        RECT 325.870 3.670 328.710 4.280 ;
        RECT 329.550 3.670 332.390 4.280 ;
        RECT 333.230 3.670 336.070 4.280 ;
        RECT 336.910 3.670 339.750 4.280 ;
        RECT 340.590 3.670 343.430 4.280 ;
        RECT 344.270 3.670 347.110 4.280 ;
        RECT 347.950 3.670 350.790 4.280 ;
        RECT 351.630 3.670 354.470 4.280 ;
        RECT 355.310 3.670 358.150 4.280 ;
        RECT 358.990 3.670 361.830 4.280 ;
        RECT 362.670 3.670 365.970 4.280 ;
        RECT 366.810 3.670 369.650 4.280 ;
        RECT 370.490 3.670 373.330 4.280 ;
        RECT 374.170 3.670 377.010 4.280 ;
        RECT 377.850 3.670 380.690 4.280 ;
        RECT 381.530 3.670 384.370 4.280 ;
        RECT 385.210 3.670 388.050 4.280 ;
        RECT 388.890 3.670 391.730 4.280 ;
        RECT 392.570 3.670 395.410 4.280 ;
        RECT 396.250 3.670 399.090 4.280 ;
        RECT 399.930 3.670 402.770 4.280 ;
        RECT 403.610 3.670 406.450 4.280 ;
        RECT 407.290 3.670 410.130 4.280 ;
        RECT 410.970 3.670 414.270 4.280 ;
        RECT 415.110 3.670 417.950 4.280 ;
        RECT 418.790 3.670 421.630 4.280 ;
        RECT 422.470 3.670 425.310 4.280 ;
        RECT 426.150 3.670 428.990 4.280 ;
        RECT 429.830 3.670 432.670 4.280 ;
        RECT 433.510 3.670 436.350 4.280 ;
        RECT 437.190 3.670 440.030 4.280 ;
        RECT 440.870 3.670 443.710 4.280 ;
        RECT 444.550 3.670 447.390 4.280 ;
        RECT 448.230 3.670 451.070 4.280 ;
        RECT 451.910 3.670 454.750 4.280 ;
        RECT 455.590 3.670 458.890 4.280 ;
        RECT 459.730 3.670 462.570 4.280 ;
        RECT 463.410 3.670 466.250 4.280 ;
        RECT 467.090 3.670 469.930 4.280 ;
        RECT 470.770 3.670 473.610 4.280 ;
        RECT 474.450 3.670 477.290 4.280 ;
        RECT 478.130 3.670 480.970 4.280 ;
        RECT 481.810 3.670 484.650 4.280 ;
        RECT 485.490 3.670 488.330 4.280 ;
        RECT 489.170 3.670 492.010 4.280 ;
        RECT 492.850 3.670 495.690 4.280 ;
        RECT 496.530 3.670 499.370 4.280 ;
        RECT 500.210 3.670 503.510 4.280 ;
        RECT 504.350 3.670 507.190 4.280 ;
        RECT 508.030 3.670 510.870 4.280 ;
        RECT 511.710 3.670 514.550 4.280 ;
        RECT 515.390 3.670 518.230 4.280 ;
        RECT 519.070 3.670 521.910 4.280 ;
        RECT 522.750 3.670 525.590 4.280 ;
        RECT 526.430 3.670 529.270 4.280 ;
        RECT 530.110 3.670 532.950 4.280 ;
        RECT 533.790 3.670 536.630 4.280 ;
        RECT 537.470 3.670 540.310 4.280 ;
        RECT 541.150 3.670 543.990 4.280 ;
        RECT 544.830 3.670 548.130 4.280 ;
        RECT 548.970 3.670 551.810 4.280 ;
        RECT 552.650 3.670 555.490 4.280 ;
        RECT 556.330 3.670 559.170 4.280 ;
        RECT 560.010 3.670 562.850 4.280 ;
        RECT 563.690 3.670 566.530 4.280 ;
        RECT 567.370 3.670 570.210 4.280 ;
        RECT 571.050 3.670 573.890 4.280 ;
        RECT 574.730 3.670 577.570 4.280 ;
        RECT 578.410 3.670 581.250 4.280 ;
        RECT 582.090 3.670 584.930 4.280 ;
        RECT 585.770 3.670 588.610 4.280 ;
        RECT 589.450 3.670 592.750 4.280 ;
        RECT 593.590 3.670 596.430 4.280 ;
        RECT 597.270 3.670 600.110 4.280 ;
        RECT 600.950 3.670 603.790 4.280 ;
        RECT 604.630 3.670 607.470 4.280 ;
        RECT 608.310 3.670 611.150 4.280 ;
        RECT 611.990 3.670 614.830 4.280 ;
        RECT 615.670 3.670 618.510 4.280 ;
        RECT 619.350 3.670 622.190 4.280 ;
        RECT 623.030 3.670 625.870 4.280 ;
        RECT 626.710 3.670 629.550 4.280 ;
        RECT 630.390 3.670 633.230 4.280 ;
        RECT 634.070 3.670 636.910 4.280 ;
        RECT 637.750 3.670 641.050 4.280 ;
        RECT 641.890 3.670 644.730 4.280 ;
        RECT 645.570 3.670 648.410 4.280 ;
        RECT 649.250 3.670 652.090 4.280 ;
        RECT 652.930 3.670 655.770 4.280 ;
        RECT 656.610 3.670 659.450 4.280 ;
        RECT 660.290 3.670 663.130 4.280 ;
        RECT 663.970 3.670 666.810 4.280 ;
        RECT 667.650 3.670 670.490 4.280 ;
        RECT 671.330 3.670 674.170 4.280 ;
        RECT 675.010 3.670 677.850 4.280 ;
        RECT 678.690 3.670 681.530 4.280 ;
        RECT 682.370 3.670 685.670 4.280 ;
        RECT 686.510 3.670 689.350 4.280 ;
        RECT 690.190 3.670 693.030 4.280 ;
        RECT 693.870 3.670 696.710 4.280 ;
        RECT 697.550 3.670 700.390 4.280 ;
        RECT 701.230 3.670 704.070 4.280 ;
        RECT 704.910 3.670 707.750 4.280 ;
        RECT 708.590 3.670 711.430 4.280 ;
        RECT 712.270 3.670 715.110 4.280 ;
        RECT 715.950 3.670 718.790 4.280 ;
        RECT 719.630 3.670 722.470 4.280 ;
        RECT 723.310 3.670 726.150 4.280 ;
        RECT 726.990 3.670 730.290 4.280 ;
        RECT 731.130 3.670 733.970 4.280 ;
        RECT 734.810 3.670 737.650 4.280 ;
        RECT 738.490 3.670 741.330 4.280 ;
        RECT 742.170 3.670 745.010 4.280 ;
        RECT 745.850 3.670 748.690 4.280 ;
        RECT 749.530 3.670 752.370 4.280 ;
        RECT 753.210 3.670 756.050 4.280 ;
        RECT 756.890 3.670 759.730 4.280 ;
        RECT 760.570 3.670 763.410 4.280 ;
        RECT 764.250 3.670 767.090 4.280 ;
        RECT 767.930 3.670 770.770 4.280 ;
        RECT 771.610 3.670 774.910 4.280 ;
        RECT 775.750 3.670 778.590 4.280 ;
        RECT 779.430 3.670 782.270 4.280 ;
        RECT 783.110 3.670 785.950 4.280 ;
        RECT 786.790 3.670 789.630 4.280 ;
        RECT 790.470 3.670 793.310 4.280 ;
        RECT 794.150 3.670 796.990 4.280 ;
        RECT 797.830 3.670 800.670 4.280 ;
        RECT 801.510 3.670 804.350 4.280 ;
        RECT 805.190 3.670 808.030 4.280 ;
        RECT 808.870 3.670 811.710 4.280 ;
        RECT 812.550 3.670 815.390 4.280 ;
        RECT 816.230 3.670 819.070 4.280 ;
        RECT 819.910 3.670 823.210 4.280 ;
        RECT 824.050 3.670 826.890 4.280 ;
        RECT 827.730 3.670 830.570 4.280 ;
        RECT 831.410 3.670 834.250 4.280 ;
        RECT 835.090 3.670 837.930 4.280 ;
        RECT 838.770 3.670 841.610 4.280 ;
        RECT 842.450 3.670 845.290 4.280 ;
        RECT 846.130 3.670 848.970 4.280 ;
        RECT 849.810 3.670 852.650 4.280 ;
        RECT 853.490 3.670 856.330 4.280 ;
        RECT 857.170 3.670 860.010 4.280 ;
        RECT 860.850 3.670 863.690 4.280 ;
        RECT 864.530 3.670 867.830 4.280 ;
        RECT 868.670 3.670 871.510 4.280 ;
        RECT 872.350 3.670 875.190 4.280 ;
        RECT 876.030 3.670 878.870 4.280 ;
        RECT 879.710 3.670 882.550 4.280 ;
        RECT 883.390 3.670 886.230 4.280 ;
        RECT 887.070 3.670 889.910 4.280 ;
        RECT 890.750 3.670 893.590 4.280 ;
        RECT 894.430 3.670 897.270 4.280 ;
        RECT 898.110 3.670 900.950 4.280 ;
        RECT 901.790 3.670 904.630 4.280 ;
        RECT 905.470 3.670 908.310 4.280 ;
        RECT 909.150 3.670 912.450 4.280 ;
        RECT 913.290 3.670 916.130 4.280 ;
        RECT 916.970 3.670 919.810 4.280 ;
        RECT 920.650 3.670 923.490 4.280 ;
        RECT 924.330 3.670 927.170 4.280 ;
        RECT 928.010 3.670 930.850 4.280 ;
        RECT 931.690 3.670 934.530 4.280 ;
        RECT 935.370 3.670 938.210 4.280 ;
        RECT 939.050 3.670 941.890 4.280 ;
        RECT 942.730 3.670 945.570 4.280 ;
        RECT 946.410 3.670 949.250 4.280 ;
        RECT 950.090 3.670 952.930 4.280 ;
        RECT 953.770 3.670 957.070 4.280 ;
        RECT 957.910 3.670 960.750 4.280 ;
        RECT 961.590 3.670 964.430 4.280 ;
        RECT 965.270 3.670 968.110 4.280 ;
        RECT 968.950 3.670 971.790 4.280 ;
        RECT 972.630 3.670 975.470 4.280 ;
        RECT 976.310 3.670 979.150 4.280 ;
        RECT 979.990 3.670 982.830 4.280 ;
        RECT 983.670 3.670 986.510 4.280 ;
        RECT 987.350 3.670 990.190 4.280 ;
        RECT 991.030 3.670 993.870 4.280 ;
        RECT 994.710 3.670 997.550 4.280 ;
      LAYER met3 ;
        RECT 4.000 1485.480 996.000 1488.005 ;
        RECT 4.000 1484.080 995.600 1485.480 ;
        RECT 4.000 1482.080 996.000 1484.080 ;
        RECT 4.400 1480.680 996.000 1482.080 ;
        RECT 4.000 1475.960 996.000 1480.680 ;
        RECT 4.000 1474.560 995.600 1475.960 ;
        RECT 4.000 1469.160 996.000 1474.560 ;
        RECT 4.400 1467.760 996.000 1469.160 ;
        RECT 4.000 1465.760 996.000 1467.760 ;
        RECT 4.000 1464.360 995.600 1465.760 ;
        RECT 4.000 1456.920 996.000 1464.360 ;
        RECT 4.400 1455.560 996.000 1456.920 ;
        RECT 4.400 1455.520 995.600 1455.560 ;
        RECT 4.000 1454.160 995.600 1455.520 ;
        RECT 4.000 1446.040 996.000 1454.160 ;
        RECT 4.000 1444.680 995.600 1446.040 ;
        RECT 4.400 1444.640 995.600 1444.680 ;
        RECT 4.400 1443.280 996.000 1444.640 ;
        RECT 4.000 1435.840 996.000 1443.280 ;
        RECT 4.000 1434.440 995.600 1435.840 ;
        RECT 4.000 1431.760 996.000 1434.440 ;
        RECT 4.400 1430.360 996.000 1431.760 ;
        RECT 4.000 1426.320 996.000 1430.360 ;
        RECT 4.000 1424.920 995.600 1426.320 ;
        RECT 4.000 1419.520 996.000 1424.920 ;
        RECT 4.400 1418.120 996.000 1419.520 ;
        RECT 4.000 1416.120 996.000 1418.120 ;
        RECT 4.000 1414.720 995.600 1416.120 ;
        RECT 4.000 1406.600 996.000 1414.720 ;
        RECT 4.400 1405.920 996.000 1406.600 ;
        RECT 4.400 1405.200 995.600 1405.920 ;
        RECT 4.000 1404.520 995.600 1405.200 ;
        RECT 4.000 1396.400 996.000 1404.520 ;
        RECT 4.000 1395.000 995.600 1396.400 ;
        RECT 4.000 1394.360 996.000 1395.000 ;
        RECT 4.400 1392.960 996.000 1394.360 ;
        RECT 4.000 1386.200 996.000 1392.960 ;
        RECT 4.000 1384.800 995.600 1386.200 ;
        RECT 4.000 1382.120 996.000 1384.800 ;
        RECT 4.400 1380.720 996.000 1382.120 ;
        RECT 4.000 1376.680 996.000 1380.720 ;
        RECT 4.000 1375.280 995.600 1376.680 ;
        RECT 4.000 1369.200 996.000 1375.280 ;
        RECT 4.400 1367.800 996.000 1369.200 ;
        RECT 4.000 1366.480 996.000 1367.800 ;
        RECT 4.000 1365.080 995.600 1366.480 ;
        RECT 4.000 1356.960 996.000 1365.080 ;
        RECT 4.400 1356.280 996.000 1356.960 ;
        RECT 4.400 1355.560 995.600 1356.280 ;
        RECT 4.000 1354.880 995.600 1355.560 ;
        RECT 4.000 1346.760 996.000 1354.880 ;
        RECT 4.000 1345.360 995.600 1346.760 ;
        RECT 4.000 1344.720 996.000 1345.360 ;
        RECT 4.400 1343.320 996.000 1344.720 ;
        RECT 4.000 1336.560 996.000 1343.320 ;
        RECT 4.000 1335.160 995.600 1336.560 ;
        RECT 4.000 1331.800 996.000 1335.160 ;
        RECT 4.400 1330.400 996.000 1331.800 ;
        RECT 4.000 1327.040 996.000 1330.400 ;
        RECT 4.000 1325.640 995.600 1327.040 ;
        RECT 4.000 1319.560 996.000 1325.640 ;
        RECT 4.400 1318.160 996.000 1319.560 ;
        RECT 4.000 1316.840 996.000 1318.160 ;
        RECT 4.000 1315.440 995.600 1316.840 ;
        RECT 4.000 1306.640 996.000 1315.440 ;
        RECT 4.400 1305.240 995.600 1306.640 ;
        RECT 4.000 1297.120 996.000 1305.240 ;
        RECT 4.000 1295.720 995.600 1297.120 ;
        RECT 4.000 1294.400 996.000 1295.720 ;
        RECT 4.400 1293.000 996.000 1294.400 ;
        RECT 4.000 1286.920 996.000 1293.000 ;
        RECT 4.000 1285.520 995.600 1286.920 ;
        RECT 4.000 1282.160 996.000 1285.520 ;
        RECT 4.400 1280.760 996.000 1282.160 ;
        RECT 4.000 1276.720 996.000 1280.760 ;
        RECT 4.000 1275.320 995.600 1276.720 ;
        RECT 4.000 1269.240 996.000 1275.320 ;
        RECT 4.400 1267.840 996.000 1269.240 ;
        RECT 4.000 1267.200 996.000 1267.840 ;
        RECT 4.000 1265.800 995.600 1267.200 ;
        RECT 4.000 1257.000 996.000 1265.800 ;
        RECT 4.400 1255.600 995.600 1257.000 ;
        RECT 4.000 1247.480 996.000 1255.600 ;
        RECT 4.000 1246.080 995.600 1247.480 ;
        RECT 4.000 1244.080 996.000 1246.080 ;
        RECT 4.400 1242.680 996.000 1244.080 ;
        RECT 4.000 1237.280 996.000 1242.680 ;
        RECT 4.000 1235.880 995.600 1237.280 ;
        RECT 4.000 1231.840 996.000 1235.880 ;
        RECT 4.400 1230.440 996.000 1231.840 ;
        RECT 4.000 1227.080 996.000 1230.440 ;
        RECT 4.000 1225.680 995.600 1227.080 ;
        RECT 4.000 1219.600 996.000 1225.680 ;
        RECT 4.400 1218.200 996.000 1219.600 ;
        RECT 4.000 1217.560 996.000 1218.200 ;
        RECT 4.000 1216.160 995.600 1217.560 ;
        RECT 4.000 1207.360 996.000 1216.160 ;
        RECT 4.000 1206.680 995.600 1207.360 ;
        RECT 4.400 1205.960 995.600 1206.680 ;
        RECT 4.400 1205.280 996.000 1205.960 ;
        RECT 4.000 1197.840 996.000 1205.280 ;
        RECT 4.000 1196.440 995.600 1197.840 ;
        RECT 4.000 1194.440 996.000 1196.440 ;
        RECT 4.400 1193.040 996.000 1194.440 ;
        RECT 4.000 1187.640 996.000 1193.040 ;
        RECT 4.000 1186.240 995.600 1187.640 ;
        RECT 4.000 1182.200 996.000 1186.240 ;
        RECT 4.400 1180.800 996.000 1182.200 ;
        RECT 4.000 1177.440 996.000 1180.800 ;
        RECT 4.000 1176.040 995.600 1177.440 ;
        RECT 4.000 1169.280 996.000 1176.040 ;
        RECT 4.400 1167.920 996.000 1169.280 ;
        RECT 4.400 1167.880 995.600 1167.920 ;
        RECT 4.000 1166.520 995.600 1167.880 ;
        RECT 4.000 1157.720 996.000 1166.520 ;
        RECT 4.000 1157.040 995.600 1157.720 ;
        RECT 4.400 1156.320 995.600 1157.040 ;
        RECT 4.400 1155.640 996.000 1156.320 ;
        RECT 4.000 1148.200 996.000 1155.640 ;
        RECT 4.000 1146.800 995.600 1148.200 ;
        RECT 4.000 1144.120 996.000 1146.800 ;
        RECT 4.400 1142.720 996.000 1144.120 ;
        RECT 4.000 1138.000 996.000 1142.720 ;
        RECT 4.000 1136.600 995.600 1138.000 ;
        RECT 4.000 1131.880 996.000 1136.600 ;
        RECT 4.400 1130.480 996.000 1131.880 ;
        RECT 4.000 1127.800 996.000 1130.480 ;
        RECT 4.000 1126.400 995.600 1127.800 ;
        RECT 4.000 1119.640 996.000 1126.400 ;
        RECT 4.400 1118.280 996.000 1119.640 ;
        RECT 4.400 1118.240 995.600 1118.280 ;
        RECT 4.000 1116.880 995.600 1118.240 ;
        RECT 4.000 1108.080 996.000 1116.880 ;
        RECT 4.000 1106.720 995.600 1108.080 ;
        RECT 4.400 1106.680 995.600 1106.720 ;
        RECT 4.400 1105.320 996.000 1106.680 ;
        RECT 4.000 1098.560 996.000 1105.320 ;
        RECT 4.000 1097.160 995.600 1098.560 ;
        RECT 4.000 1094.480 996.000 1097.160 ;
        RECT 4.400 1093.080 996.000 1094.480 ;
        RECT 4.000 1088.360 996.000 1093.080 ;
        RECT 4.000 1086.960 995.600 1088.360 ;
        RECT 4.000 1081.560 996.000 1086.960 ;
        RECT 4.400 1080.160 996.000 1081.560 ;
        RECT 4.000 1078.160 996.000 1080.160 ;
        RECT 4.000 1076.760 995.600 1078.160 ;
        RECT 4.000 1069.320 996.000 1076.760 ;
        RECT 4.400 1068.640 996.000 1069.320 ;
        RECT 4.400 1067.920 995.600 1068.640 ;
        RECT 4.000 1067.240 995.600 1067.920 ;
        RECT 4.000 1058.440 996.000 1067.240 ;
        RECT 4.000 1057.080 995.600 1058.440 ;
        RECT 4.400 1057.040 995.600 1057.080 ;
        RECT 4.400 1055.680 996.000 1057.040 ;
        RECT 4.000 1048.240 996.000 1055.680 ;
        RECT 4.000 1046.840 995.600 1048.240 ;
        RECT 4.000 1044.160 996.000 1046.840 ;
        RECT 4.400 1042.760 996.000 1044.160 ;
        RECT 4.000 1038.720 996.000 1042.760 ;
        RECT 4.000 1037.320 995.600 1038.720 ;
        RECT 4.000 1031.920 996.000 1037.320 ;
        RECT 4.400 1030.520 996.000 1031.920 ;
        RECT 4.000 1028.520 996.000 1030.520 ;
        RECT 4.000 1027.120 995.600 1028.520 ;
        RECT 4.000 1019.680 996.000 1027.120 ;
        RECT 4.400 1019.000 996.000 1019.680 ;
        RECT 4.400 1018.280 995.600 1019.000 ;
        RECT 4.000 1017.600 995.600 1018.280 ;
        RECT 4.000 1008.800 996.000 1017.600 ;
        RECT 4.000 1007.400 995.600 1008.800 ;
        RECT 4.000 1006.760 996.000 1007.400 ;
        RECT 4.400 1005.360 996.000 1006.760 ;
        RECT 4.000 998.600 996.000 1005.360 ;
        RECT 4.000 997.200 995.600 998.600 ;
        RECT 4.000 994.520 996.000 997.200 ;
        RECT 4.400 993.120 996.000 994.520 ;
        RECT 4.000 989.080 996.000 993.120 ;
        RECT 4.000 987.680 995.600 989.080 ;
        RECT 4.000 981.600 996.000 987.680 ;
        RECT 4.400 980.200 996.000 981.600 ;
        RECT 4.000 978.880 996.000 980.200 ;
        RECT 4.000 977.480 995.600 978.880 ;
        RECT 4.000 969.360 996.000 977.480 ;
        RECT 4.400 967.960 995.600 969.360 ;
        RECT 4.000 959.160 996.000 967.960 ;
        RECT 4.000 957.760 995.600 959.160 ;
        RECT 4.000 957.120 996.000 957.760 ;
        RECT 4.400 955.720 996.000 957.120 ;
        RECT 4.000 948.960 996.000 955.720 ;
        RECT 4.000 947.560 995.600 948.960 ;
        RECT 4.000 944.200 996.000 947.560 ;
        RECT 4.400 942.800 996.000 944.200 ;
        RECT 4.000 939.440 996.000 942.800 ;
        RECT 4.000 938.040 995.600 939.440 ;
        RECT 4.000 931.960 996.000 938.040 ;
        RECT 4.400 930.560 996.000 931.960 ;
        RECT 4.000 929.240 996.000 930.560 ;
        RECT 4.000 927.840 995.600 929.240 ;
        RECT 4.000 919.720 996.000 927.840 ;
        RECT 4.000 919.040 995.600 919.720 ;
        RECT 4.400 918.320 995.600 919.040 ;
        RECT 4.400 917.640 996.000 918.320 ;
        RECT 4.000 909.520 996.000 917.640 ;
        RECT 4.000 908.120 995.600 909.520 ;
        RECT 4.000 906.800 996.000 908.120 ;
        RECT 4.400 905.400 996.000 906.800 ;
        RECT 4.000 899.320 996.000 905.400 ;
        RECT 4.000 897.920 995.600 899.320 ;
        RECT 4.000 894.560 996.000 897.920 ;
        RECT 4.400 893.160 996.000 894.560 ;
        RECT 4.000 889.800 996.000 893.160 ;
        RECT 4.000 888.400 995.600 889.800 ;
        RECT 4.000 881.640 996.000 888.400 ;
        RECT 4.400 880.240 996.000 881.640 ;
        RECT 4.000 879.600 996.000 880.240 ;
        RECT 4.000 878.200 995.600 879.600 ;
        RECT 4.000 870.080 996.000 878.200 ;
        RECT 4.000 869.400 995.600 870.080 ;
        RECT 4.400 868.680 995.600 869.400 ;
        RECT 4.400 868.000 996.000 868.680 ;
        RECT 4.000 859.880 996.000 868.000 ;
        RECT 4.000 858.480 995.600 859.880 ;
        RECT 4.000 857.160 996.000 858.480 ;
        RECT 4.400 855.760 996.000 857.160 ;
        RECT 4.000 849.680 996.000 855.760 ;
        RECT 4.000 848.280 995.600 849.680 ;
        RECT 4.000 844.240 996.000 848.280 ;
        RECT 4.400 842.840 996.000 844.240 ;
        RECT 4.000 840.160 996.000 842.840 ;
        RECT 4.000 838.760 995.600 840.160 ;
        RECT 4.000 832.000 996.000 838.760 ;
        RECT 4.400 830.600 996.000 832.000 ;
        RECT 4.000 829.960 996.000 830.600 ;
        RECT 4.000 828.560 995.600 829.960 ;
        RECT 4.000 819.760 996.000 828.560 ;
        RECT 4.000 819.080 995.600 819.760 ;
        RECT 4.400 818.360 995.600 819.080 ;
        RECT 4.400 817.680 996.000 818.360 ;
        RECT 4.000 810.240 996.000 817.680 ;
        RECT 4.000 808.840 995.600 810.240 ;
        RECT 4.000 806.840 996.000 808.840 ;
        RECT 4.400 805.440 996.000 806.840 ;
        RECT 4.000 800.040 996.000 805.440 ;
        RECT 4.000 798.640 995.600 800.040 ;
        RECT 4.000 794.600 996.000 798.640 ;
        RECT 4.400 793.200 996.000 794.600 ;
        RECT 4.000 790.520 996.000 793.200 ;
        RECT 4.000 789.120 995.600 790.520 ;
        RECT 4.000 781.680 996.000 789.120 ;
        RECT 4.400 780.320 996.000 781.680 ;
        RECT 4.400 780.280 995.600 780.320 ;
        RECT 4.000 778.920 995.600 780.280 ;
        RECT 4.000 770.120 996.000 778.920 ;
        RECT 4.000 769.440 995.600 770.120 ;
        RECT 4.400 768.720 995.600 769.440 ;
        RECT 4.400 768.040 996.000 768.720 ;
        RECT 4.000 760.600 996.000 768.040 ;
        RECT 4.000 759.200 995.600 760.600 ;
        RECT 4.000 757.200 996.000 759.200 ;
        RECT 4.400 755.800 996.000 757.200 ;
        RECT 4.000 750.400 996.000 755.800 ;
        RECT 4.000 749.000 995.600 750.400 ;
        RECT 4.000 744.280 996.000 749.000 ;
        RECT 4.400 742.880 996.000 744.280 ;
        RECT 4.000 740.880 996.000 742.880 ;
        RECT 4.000 739.480 995.600 740.880 ;
        RECT 4.000 732.040 996.000 739.480 ;
        RECT 4.400 730.680 996.000 732.040 ;
        RECT 4.400 730.640 995.600 730.680 ;
        RECT 4.000 729.280 995.600 730.640 ;
        RECT 4.000 720.480 996.000 729.280 ;
        RECT 4.000 719.120 995.600 720.480 ;
        RECT 4.400 719.080 995.600 719.120 ;
        RECT 4.400 717.720 996.000 719.080 ;
        RECT 4.000 710.960 996.000 717.720 ;
        RECT 4.000 709.560 995.600 710.960 ;
        RECT 4.000 706.880 996.000 709.560 ;
        RECT 4.400 705.480 996.000 706.880 ;
        RECT 4.000 700.760 996.000 705.480 ;
        RECT 4.000 699.360 995.600 700.760 ;
        RECT 4.000 694.640 996.000 699.360 ;
        RECT 4.400 693.240 996.000 694.640 ;
        RECT 4.000 691.240 996.000 693.240 ;
        RECT 4.000 689.840 995.600 691.240 ;
        RECT 4.000 681.720 996.000 689.840 ;
        RECT 4.400 681.040 996.000 681.720 ;
        RECT 4.400 680.320 995.600 681.040 ;
        RECT 4.000 679.640 995.600 680.320 ;
        RECT 4.000 670.840 996.000 679.640 ;
        RECT 4.000 669.480 995.600 670.840 ;
        RECT 4.400 669.440 995.600 669.480 ;
        RECT 4.400 668.080 996.000 669.440 ;
        RECT 4.000 661.320 996.000 668.080 ;
        RECT 4.000 659.920 995.600 661.320 ;
        RECT 4.000 656.560 996.000 659.920 ;
        RECT 4.400 655.160 996.000 656.560 ;
        RECT 4.000 651.120 996.000 655.160 ;
        RECT 4.000 649.720 995.600 651.120 ;
        RECT 4.000 644.320 996.000 649.720 ;
        RECT 4.400 642.920 996.000 644.320 ;
        RECT 4.000 640.920 996.000 642.920 ;
        RECT 4.000 639.520 995.600 640.920 ;
        RECT 4.000 632.080 996.000 639.520 ;
        RECT 4.400 631.400 996.000 632.080 ;
        RECT 4.400 630.680 995.600 631.400 ;
        RECT 4.000 630.000 995.600 630.680 ;
        RECT 4.000 621.200 996.000 630.000 ;
        RECT 4.000 619.800 995.600 621.200 ;
        RECT 4.000 619.160 996.000 619.800 ;
        RECT 4.400 617.760 996.000 619.160 ;
        RECT 4.000 611.680 996.000 617.760 ;
        RECT 4.000 610.280 995.600 611.680 ;
        RECT 4.000 606.920 996.000 610.280 ;
        RECT 4.400 605.520 996.000 606.920 ;
        RECT 4.000 601.480 996.000 605.520 ;
        RECT 4.000 600.080 995.600 601.480 ;
        RECT 4.000 594.680 996.000 600.080 ;
        RECT 4.400 593.280 996.000 594.680 ;
        RECT 4.000 591.280 996.000 593.280 ;
        RECT 4.000 589.880 995.600 591.280 ;
        RECT 4.000 581.760 996.000 589.880 ;
        RECT 4.400 580.360 995.600 581.760 ;
        RECT 4.000 571.560 996.000 580.360 ;
        RECT 4.000 570.160 995.600 571.560 ;
        RECT 4.000 569.520 996.000 570.160 ;
        RECT 4.400 568.120 996.000 569.520 ;
        RECT 4.000 562.040 996.000 568.120 ;
        RECT 4.000 560.640 995.600 562.040 ;
        RECT 4.000 556.600 996.000 560.640 ;
        RECT 4.400 555.200 996.000 556.600 ;
        RECT 4.000 551.840 996.000 555.200 ;
        RECT 4.000 550.440 995.600 551.840 ;
        RECT 4.000 544.360 996.000 550.440 ;
        RECT 4.400 542.960 996.000 544.360 ;
        RECT 4.000 541.640 996.000 542.960 ;
        RECT 4.000 540.240 995.600 541.640 ;
        RECT 4.000 532.120 996.000 540.240 ;
        RECT 4.400 530.720 995.600 532.120 ;
        RECT 4.000 521.920 996.000 530.720 ;
        RECT 4.000 520.520 995.600 521.920 ;
        RECT 4.000 519.200 996.000 520.520 ;
        RECT 4.400 517.800 996.000 519.200 ;
        RECT 4.000 512.400 996.000 517.800 ;
        RECT 4.000 511.000 995.600 512.400 ;
        RECT 4.000 506.960 996.000 511.000 ;
        RECT 4.400 505.560 996.000 506.960 ;
        RECT 4.000 502.200 996.000 505.560 ;
        RECT 4.000 500.800 995.600 502.200 ;
        RECT 4.000 494.040 996.000 500.800 ;
        RECT 4.400 492.640 996.000 494.040 ;
        RECT 4.000 492.000 996.000 492.640 ;
        RECT 4.000 490.600 995.600 492.000 ;
        RECT 4.000 482.480 996.000 490.600 ;
        RECT 4.000 481.800 995.600 482.480 ;
        RECT 4.400 481.080 995.600 481.800 ;
        RECT 4.400 480.400 996.000 481.080 ;
        RECT 4.000 472.280 996.000 480.400 ;
        RECT 4.000 470.880 995.600 472.280 ;
        RECT 4.000 469.560 996.000 470.880 ;
        RECT 4.400 468.160 996.000 469.560 ;
        RECT 4.000 462.760 996.000 468.160 ;
        RECT 4.000 461.360 995.600 462.760 ;
        RECT 4.000 456.640 996.000 461.360 ;
        RECT 4.400 455.240 996.000 456.640 ;
        RECT 4.000 452.560 996.000 455.240 ;
        RECT 4.000 451.160 995.600 452.560 ;
        RECT 4.000 444.400 996.000 451.160 ;
        RECT 4.400 443.000 996.000 444.400 ;
        RECT 4.000 442.360 996.000 443.000 ;
        RECT 4.000 440.960 995.600 442.360 ;
        RECT 4.000 432.840 996.000 440.960 ;
        RECT 4.000 432.160 995.600 432.840 ;
        RECT 4.400 431.440 995.600 432.160 ;
        RECT 4.400 430.760 996.000 431.440 ;
        RECT 4.000 422.640 996.000 430.760 ;
        RECT 4.000 421.240 995.600 422.640 ;
        RECT 4.000 419.240 996.000 421.240 ;
        RECT 4.400 417.840 996.000 419.240 ;
        RECT 4.000 412.440 996.000 417.840 ;
        RECT 4.000 411.040 995.600 412.440 ;
        RECT 4.000 407.000 996.000 411.040 ;
        RECT 4.400 405.600 996.000 407.000 ;
        RECT 4.000 402.920 996.000 405.600 ;
        RECT 4.000 401.520 995.600 402.920 ;
        RECT 4.000 394.080 996.000 401.520 ;
        RECT 4.400 392.720 996.000 394.080 ;
        RECT 4.400 392.680 995.600 392.720 ;
        RECT 4.000 391.320 995.600 392.680 ;
        RECT 4.000 383.200 996.000 391.320 ;
        RECT 4.000 381.840 995.600 383.200 ;
        RECT 4.400 381.800 995.600 381.840 ;
        RECT 4.400 380.440 996.000 381.800 ;
        RECT 4.000 373.000 996.000 380.440 ;
        RECT 4.000 371.600 995.600 373.000 ;
        RECT 4.000 369.600 996.000 371.600 ;
        RECT 4.400 368.200 996.000 369.600 ;
        RECT 4.000 362.800 996.000 368.200 ;
        RECT 4.000 361.400 995.600 362.800 ;
        RECT 4.000 356.680 996.000 361.400 ;
        RECT 4.400 355.280 996.000 356.680 ;
        RECT 4.000 353.280 996.000 355.280 ;
        RECT 4.000 351.880 995.600 353.280 ;
        RECT 4.000 344.440 996.000 351.880 ;
        RECT 4.400 343.080 996.000 344.440 ;
        RECT 4.400 343.040 995.600 343.080 ;
        RECT 4.000 341.680 995.600 343.040 ;
        RECT 4.000 333.560 996.000 341.680 ;
        RECT 4.000 332.160 995.600 333.560 ;
        RECT 4.000 331.520 996.000 332.160 ;
        RECT 4.400 330.120 996.000 331.520 ;
        RECT 4.000 323.360 996.000 330.120 ;
        RECT 4.000 321.960 995.600 323.360 ;
        RECT 4.000 319.280 996.000 321.960 ;
        RECT 4.400 317.880 996.000 319.280 ;
        RECT 4.000 313.160 996.000 317.880 ;
        RECT 4.000 311.760 995.600 313.160 ;
        RECT 4.000 307.040 996.000 311.760 ;
        RECT 4.400 305.640 996.000 307.040 ;
        RECT 4.000 303.640 996.000 305.640 ;
        RECT 4.000 302.240 995.600 303.640 ;
        RECT 4.000 294.120 996.000 302.240 ;
        RECT 4.400 293.440 996.000 294.120 ;
        RECT 4.400 292.720 995.600 293.440 ;
        RECT 4.000 292.040 995.600 292.720 ;
        RECT 4.000 283.920 996.000 292.040 ;
        RECT 4.000 282.520 995.600 283.920 ;
        RECT 4.000 281.880 996.000 282.520 ;
        RECT 4.400 280.480 996.000 281.880 ;
        RECT 4.000 273.720 996.000 280.480 ;
        RECT 4.000 272.320 995.600 273.720 ;
        RECT 4.000 269.640 996.000 272.320 ;
        RECT 4.400 268.240 996.000 269.640 ;
        RECT 4.000 263.520 996.000 268.240 ;
        RECT 4.000 262.120 995.600 263.520 ;
        RECT 4.000 256.720 996.000 262.120 ;
        RECT 4.400 255.320 996.000 256.720 ;
        RECT 4.000 254.000 996.000 255.320 ;
        RECT 4.000 252.600 995.600 254.000 ;
        RECT 4.000 244.480 996.000 252.600 ;
        RECT 4.400 243.800 996.000 244.480 ;
        RECT 4.400 243.080 995.600 243.800 ;
        RECT 4.000 242.400 995.600 243.080 ;
        RECT 4.000 234.280 996.000 242.400 ;
        RECT 4.000 232.880 995.600 234.280 ;
        RECT 4.000 231.560 996.000 232.880 ;
        RECT 4.400 230.160 996.000 231.560 ;
        RECT 4.000 224.080 996.000 230.160 ;
        RECT 4.000 222.680 995.600 224.080 ;
        RECT 4.000 219.320 996.000 222.680 ;
        RECT 4.400 217.920 996.000 219.320 ;
        RECT 4.000 213.880 996.000 217.920 ;
        RECT 4.000 212.480 995.600 213.880 ;
        RECT 4.000 207.080 996.000 212.480 ;
        RECT 4.400 205.680 996.000 207.080 ;
        RECT 4.000 204.360 996.000 205.680 ;
        RECT 4.000 202.960 995.600 204.360 ;
        RECT 4.000 194.160 996.000 202.960 ;
        RECT 4.400 192.760 995.600 194.160 ;
        RECT 4.000 183.960 996.000 192.760 ;
        RECT 4.000 182.560 995.600 183.960 ;
        RECT 4.000 181.920 996.000 182.560 ;
        RECT 4.400 180.520 996.000 181.920 ;
        RECT 4.000 174.440 996.000 180.520 ;
        RECT 4.000 173.040 995.600 174.440 ;
        RECT 4.000 169.000 996.000 173.040 ;
        RECT 4.400 167.600 996.000 169.000 ;
        RECT 4.000 164.240 996.000 167.600 ;
        RECT 4.000 162.840 995.600 164.240 ;
        RECT 4.000 156.760 996.000 162.840 ;
        RECT 4.400 155.360 996.000 156.760 ;
        RECT 4.000 154.720 996.000 155.360 ;
        RECT 4.000 153.320 995.600 154.720 ;
        RECT 4.000 144.520 996.000 153.320 ;
        RECT 4.400 143.120 995.600 144.520 ;
        RECT 4.000 134.320 996.000 143.120 ;
        RECT 4.000 132.920 995.600 134.320 ;
        RECT 4.000 131.600 996.000 132.920 ;
        RECT 4.400 130.200 996.000 131.600 ;
        RECT 4.000 124.800 996.000 130.200 ;
        RECT 4.000 123.400 995.600 124.800 ;
        RECT 4.000 119.360 996.000 123.400 ;
        RECT 4.400 117.960 996.000 119.360 ;
        RECT 4.000 114.600 996.000 117.960 ;
        RECT 4.000 113.200 995.600 114.600 ;
        RECT 4.000 107.120 996.000 113.200 ;
        RECT 4.400 105.720 996.000 107.120 ;
        RECT 4.000 105.080 996.000 105.720 ;
        RECT 4.000 103.680 995.600 105.080 ;
        RECT 4.000 94.880 996.000 103.680 ;
        RECT 4.000 94.200 995.600 94.880 ;
        RECT 4.400 93.480 995.600 94.200 ;
        RECT 4.400 92.800 996.000 93.480 ;
        RECT 4.000 84.680 996.000 92.800 ;
        RECT 4.000 83.280 995.600 84.680 ;
        RECT 4.000 81.960 996.000 83.280 ;
        RECT 4.400 80.560 996.000 81.960 ;
        RECT 4.000 75.160 996.000 80.560 ;
        RECT 4.000 73.760 995.600 75.160 ;
        RECT 4.000 69.040 996.000 73.760 ;
        RECT 4.400 67.640 996.000 69.040 ;
        RECT 4.000 64.960 996.000 67.640 ;
        RECT 4.000 63.560 995.600 64.960 ;
        RECT 4.000 56.800 996.000 63.560 ;
        RECT 4.400 55.440 996.000 56.800 ;
        RECT 4.400 55.400 995.600 55.440 ;
        RECT 4.000 54.040 995.600 55.400 ;
        RECT 4.000 45.240 996.000 54.040 ;
        RECT 4.000 44.560 995.600 45.240 ;
        RECT 4.400 43.840 995.600 44.560 ;
        RECT 4.400 43.160 996.000 43.840 ;
        RECT 4.000 35.040 996.000 43.160 ;
        RECT 4.000 33.640 995.600 35.040 ;
        RECT 4.000 31.640 996.000 33.640 ;
        RECT 4.400 30.240 996.000 31.640 ;
        RECT 4.000 25.520 996.000 30.240 ;
        RECT 4.000 24.120 995.600 25.520 ;
        RECT 4.000 19.400 996.000 24.120 ;
        RECT 4.400 18.000 996.000 19.400 ;
        RECT 4.000 15.320 996.000 18.000 ;
        RECT 4.000 13.920 995.600 15.320 ;
        RECT 4.000 7.160 996.000 13.920 ;
        RECT 4.400 6.295 996.000 7.160 ;
      LAYER met4 ;
        RECT 303.895 10.240 327.840 214.705 ;
        RECT 330.240 10.240 404.640 214.705 ;
        RECT 407.040 10.240 481.440 214.705 ;
        RECT 483.840 10.240 558.240 214.705 ;
        RECT 560.640 10.240 565.505 214.705 ;
        RECT 303.895 6.295 565.505 10.240 ;
  END
END user_proj_example
END LIBRARY

