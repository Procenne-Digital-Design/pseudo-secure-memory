magic
tech sky130A
magscale 1 2
timestamp 1647413277
<< viali >>
rect 4629 117317 4663 117351
rect 1869 117249 1903 117283
rect 7849 117249 7883 117283
rect 11713 117249 11747 117283
rect 15577 117249 15611 117283
rect 19441 117249 19475 117283
rect 22661 117249 22695 117283
rect 27169 117249 27203 117283
rect 30389 117249 30423 117283
rect 34713 117249 34747 117283
rect 35265 117249 35299 117283
rect 37473 117249 37507 117283
rect 41337 117249 41371 117283
rect 45201 117249 45235 117283
rect 49249 117249 49283 117283
rect 52745 117249 52779 117283
rect 56149 117249 56183 117283
rect 60657 117249 60691 117283
rect 63877 117249 63911 117283
rect 67097 117249 67131 117283
rect 71237 117249 71271 117283
rect 74825 117249 74859 117283
rect 77125 117249 77159 117283
rect 5457 117181 5491 117215
rect 11897 117181 11931 117215
rect 56333 117181 56367 117215
rect 77401 117181 77435 117215
rect 19625 117113 19659 117147
rect 22845 117113 22879 117147
rect 30573 117113 30607 117147
rect 34897 117113 34931 117147
rect 37657 117113 37691 117147
rect 45385 117113 45419 117147
rect 52929 117113 52963 117147
rect 60473 117113 60507 117147
rect 67281 117113 67315 117147
rect 75009 117113 75043 117147
rect 2145 117045 2179 117079
rect 8033 117045 8067 117079
rect 15761 117045 15795 117079
rect 26985 117045 27019 117079
rect 41521 117045 41555 117079
rect 49065 117045 49099 117079
rect 64061 117045 64095 117079
rect 66729 117045 66763 117079
rect 71329 117045 71363 117079
rect 74549 117045 74583 117079
rect 78045 116841 78079 116875
rect 1869 116637 1903 116671
rect 77861 116637 77895 116671
rect 2237 116569 2271 116603
rect 40785 116297 40819 116331
rect 39865 116161 39899 116195
rect 40693 116161 40727 116195
rect 40049 116025 40083 116059
rect 77861 114461 77895 114495
rect 78045 114325 78079 114359
rect 24225 114121 24259 114155
rect 24409 113985 24443 114019
rect 1409 113373 1443 113407
rect 1593 113237 1627 113271
rect 66545 111877 66579 111911
rect 66729 111809 66763 111843
rect 77677 110721 77711 110755
rect 77861 110517 77895 110551
rect 1869 109633 1903 109667
rect 1961 109429 1995 109463
rect 40049 109225 40083 109259
rect 39865 109021 39899 109055
rect 77677 106369 77711 106403
rect 77861 106165 77895 106199
rect 1409 105757 1443 105791
rect 1685 105689 1719 105723
rect 77861 103717 77895 103751
rect 78045 103581 78079 103615
rect 77677 103105 77711 103139
rect 77309 102901 77343 102935
rect 77861 102901 77895 102935
rect 1409 101405 1443 101439
rect 1593 101269 1627 101303
rect 58633 100521 58667 100555
rect 58541 100249 58575 100283
rect 77677 98753 77711 98787
rect 77861 98617 77895 98651
rect 1409 97665 1443 97699
rect 1685 97597 1719 97631
rect 40325 95897 40359 95931
rect 40417 95829 40451 95863
rect 77861 94877 77895 94911
rect 78045 94741 78079 94775
rect 1409 94401 1443 94435
rect 1593 94197 1627 94231
rect 41429 92361 41463 92395
rect 41337 92225 41371 92259
rect 77953 90457 77987 90491
rect 78045 90389 78079 90423
rect 1501 90049 1535 90083
rect 2053 89981 2087 90015
rect 39957 88961 39991 88995
rect 40049 88757 40083 88791
rect 77769 87193 77803 87227
rect 77861 87125 77895 87159
rect 1409 86173 1443 86207
rect 1593 86037 1627 86071
rect 77677 83521 77711 83555
rect 77861 83317 77895 83351
rect 1409 81821 1443 81855
rect 1685 81753 1719 81787
rect 10701 79305 10735 79339
rect 10609 79169 10643 79203
rect 77585 79169 77619 79203
rect 77677 78965 77711 78999
rect 1409 78557 1443 78591
rect 1593 78421 1627 78455
rect 2605 78217 2639 78251
rect 2789 78081 2823 78115
rect 77861 75293 77895 75327
rect 78045 75157 78079 75191
rect 1409 74205 1443 74239
rect 1593 74069 1627 74103
rect 67833 72029 67867 72063
rect 68109 71961 68143 71995
rect 77677 71553 77711 71587
rect 77861 71417 77895 71451
rect 76573 71145 76607 71179
rect 2053 71077 2087 71111
rect 76757 70941 76791 70975
rect 1869 70873 1903 70907
rect 1409 70465 1443 70499
rect 1593 70261 1627 70295
rect 1777 70057 1811 70091
rect 1961 69853 1995 69887
rect 77769 67609 77803 67643
rect 77861 67541 77895 67575
rect 1409 66113 1443 66147
rect 2329 66113 2363 66147
rect 1593 65977 1627 66011
rect 2145 65977 2179 66011
rect 41889 65569 41923 65603
rect 1869 65501 1903 65535
rect 39865 65501 39899 65535
rect 40141 65433 40175 65467
rect 1961 65365 1995 65399
rect 40049 65161 40083 65195
rect 41061 65161 41095 65195
rect 40233 65025 40267 65059
rect 40693 64957 40727 64991
rect 41245 64889 41279 64923
rect 41061 64821 41095 64855
rect 40049 64413 40083 64447
rect 40509 64413 40543 64447
rect 40785 64413 40819 64447
rect 40877 64413 40911 64447
rect 39497 63937 39531 63971
rect 39589 63733 39623 63767
rect 77493 63325 77527 63359
rect 77861 63325 77895 63359
rect 78045 63189 78079 63223
rect 1409 62849 1443 62883
rect 1593 62645 1627 62679
rect 39865 61149 39899 61183
rect 40141 61081 40175 61115
rect 39957 60741 39991 60775
rect 40877 60741 40911 60775
rect 38945 60673 38979 60707
rect 39221 60605 39255 60639
rect 40141 60537 40175 60571
rect 41153 60469 41187 60503
rect 35817 60265 35851 60299
rect 36369 60265 36403 60299
rect 38301 60265 38335 60299
rect 77861 60265 77895 60299
rect 41245 60129 41279 60163
rect 1777 60061 1811 60095
rect 19257 60061 19291 60095
rect 38117 60061 38151 60095
rect 39957 60061 39991 60095
rect 41061 60061 41095 60095
rect 62957 60061 62991 60095
rect 19533 59993 19567 60027
rect 35173 59993 35207 60027
rect 36277 59993 36311 60027
rect 38945 59993 38979 60027
rect 40509 59993 40543 60027
rect 77769 59993 77803 60027
rect 1961 59925 1995 59959
rect 35265 59925 35299 59959
rect 37749 59925 37783 59959
rect 39221 59925 39255 59959
rect 63049 59925 63083 59959
rect 77769 59721 77803 59755
rect 38669 59585 38703 59619
rect 38945 59585 38979 59619
rect 39957 59585 39991 59619
rect 41061 59585 41095 59619
rect 74733 59585 74767 59619
rect 77953 59585 77987 59619
rect 39129 59517 39163 59551
rect 40509 59517 40543 59551
rect 41245 59449 41279 59483
rect 74549 59381 74583 59415
rect 2973 59177 3007 59211
rect 1409 58973 1443 59007
rect 2789 58973 2823 59007
rect 39865 58973 39899 59007
rect 40141 58905 40175 58939
rect 1593 58837 1627 58871
rect 2789 58633 2823 58667
rect 2973 58497 3007 58531
rect 77677 56321 77711 56355
rect 77861 56117 77895 56151
rect 1685 54621 1719 54655
rect 2053 54621 2087 54655
rect 1501 54485 1535 54519
rect 77677 51969 77711 52003
rect 77861 51765 77895 51799
rect 1685 50881 1719 50915
rect 2053 50881 2087 50915
rect 1501 50677 1535 50711
rect 1593 47141 1627 47175
rect 1409 47005 1443 47039
rect 77861 43741 77895 43775
rect 78045 43605 78079 43639
rect 1869 43265 1903 43299
rect 2145 43061 2179 43095
rect 77769 42721 77803 42755
rect 77585 42585 77619 42619
rect 77861 40477 77895 40511
rect 78045 40341 78079 40375
rect 77493 40137 77527 40171
rect 77677 40001 77711 40035
rect 1869 38913 1903 38947
rect 2145 38709 2179 38743
rect 77861 36125 77895 36159
rect 78045 35989 78079 36023
rect 1409 35037 1443 35071
rect 1593 34901 1627 34935
rect 71881 34629 71915 34663
rect 71697 34561 71731 34595
rect 77861 33065 77895 33099
rect 78045 32861 78079 32895
rect 77677 32385 77711 32419
rect 77861 32181 77895 32215
rect 1685 31841 1719 31875
rect 1409 31773 1443 31807
rect 77769 28169 77803 28203
rect 77953 28033 77987 28067
rect 1409 27421 1443 27455
rect 1685 27353 1719 27387
rect 39589 25857 39623 25891
rect 40233 25857 40267 25891
rect 39957 25653 39991 25687
rect 77677 24769 77711 24803
rect 77309 24565 77343 24599
rect 77861 24565 77895 24599
rect 1409 23681 1443 23715
rect 1685 23613 1719 23647
rect 77861 20893 77895 20927
rect 78045 20757 78079 20791
rect 1409 19329 1443 19363
rect 1593 19125 1627 19159
rect 77861 16541 77895 16575
rect 78045 16405 78079 16439
rect 1961 16201 1995 16235
rect 1685 16065 1719 16099
rect 1501 15861 1535 15895
rect 2881 13481 2915 13515
rect 2697 13277 2731 13311
rect 77769 12869 77803 12903
rect 77493 12801 77527 12835
rect 40325 12121 40359 12155
rect 40601 12053 40635 12087
rect 1685 11781 1719 11815
rect 1409 11713 1443 11747
rect 78045 10081 78079 10115
rect 77493 10013 77527 10047
rect 77861 8925 77895 8959
rect 77493 8789 77527 8823
rect 78045 8789 78079 8823
rect 1409 7837 1443 7871
rect 1593 7701 1627 7735
rect 2421 7497 2455 7531
rect 2697 7497 2731 7531
rect 2881 7361 2915 7395
rect 77677 5185 77711 5219
rect 77861 4981 77895 5015
rect 77861 4777 77895 4811
rect 78045 4573 78079 4607
rect 1685 3553 1719 3587
rect 1409 3485 1443 3519
rect 15117 3485 15151 3519
rect 40969 3485 41003 3519
rect 41889 3485 41923 3519
rect 40325 3417 40359 3451
rect 14933 3349 14967 3383
rect 40417 3349 40451 3383
rect 41153 3349 41187 3383
rect 41705 3349 41739 3383
rect 77309 3009 77343 3043
rect 77585 2941 77619 2975
rect 18337 2601 18371 2635
rect 29929 2601 29963 2635
rect 33149 2601 33183 2635
rect 47777 2601 47811 2635
rect 66637 2601 66671 2635
rect 15209 2533 15243 2567
rect 1685 2465 1719 2499
rect 4445 2465 4479 2499
rect 71145 2465 71179 2499
rect 77401 2465 77435 2499
rect 1409 2397 1443 2431
rect 3893 2397 3927 2431
rect 7297 2397 7331 2431
rect 11529 2397 11563 2431
rect 22017 2397 22051 2431
rect 25881 2397 25915 2431
rect 29745 2397 29779 2431
rect 37289 2397 37323 2431
rect 40693 2397 40727 2431
rect 45017 2397 45051 2431
rect 47961 2397 47995 2431
rect 51641 2397 51675 2431
rect 55505 2397 55539 2431
rect 55781 2397 55815 2431
rect 59093 2397 59127 2431
rect 59369 2397 59403 2431
rect 63049 2397 63083 2431
rect 66453 2397 66487 2431
rect 70869 2397 70903 2431
rect 73813 2397 73847 2431
rect 74181 2397 74215 2431
rect 77125 2397 77159 2431
rect 7849 2329 7883 2363
rect 15025 2329 15059 2363
rect 18245 2329 18279 2363
rect 33057 2329 33091 2363
rect 45293 2329 45327 2363
rect 51917 2329 51951 2363
rect 63877 2329 63911 2363
rect 11713 2261 11747 2295
rect 22201 2261 22235 2295
rect 26065 2261 26099 2295
rect 37473 2261 37507 2295
rect 40877 2261 40911 2295
rect 74365 2261 74399 2295
<< metal1 >>
rect 1104 117530 78844 117552
rect 1104 117478 19574 117530
rect 19626 117478 19638 117530
rect 19690 117478 19702 117530
rect 19754 117478 19766 117530
rect 19818 117478 19830 117530
rect 19882 117478 50294 117530
rect 50346 117478 50358 117530
rect 50410 117478 50422 117530
rect 50474 117478 50486 117530
rect 50538 117478 50550 117530
rect 50602 117478 78844 117530
rect 1104 117456 78844 117478
rect 4614 117348 4620 117360
rect 4575 117320 4620 117348
rect 4614 117308 4620 117320
rect 4672 117308 4678 117360
rect 658 117240 664 117292
rect 716 117280 722 117292
rect 1857 117283 1915 117289
rect 1857 117280 1869 117283
rect 716 117252 1869 117280
rect 716 117240 722 117252
rect 1857 117249 1869 117252
rect 1903 117249 1915 117283
rect 7834 117280 7840 117292
rect 7795 117252 7840 117280
rect 1857 117243 1915 117249
rect 7834 117240 7840 117252
rect 7892 117240 7898 117292
rect 11698 117280 11704 117292
rect 11659 117252 11704 117280
rect 11698 117240 11704 117252
rect 11756 117240 11762 117292
rect 15562 117280 15568 117292
rect 15523 117252 15568 117280
rect 15562 117240 15568 117252
rect 15620 117240 15626 117292
rect 19426 117280 19432 117292
rect 19387 117252 19432 117280
rect 19426 117240 19432 117252
rect 19484 117240 19490 117292
rect 22646 117280 22652 117292
rect 22607 117252 22652 117280
rect 22646 117240 22652 117252
rect 22704 117240 22710 117292
rect 26418 117240 26424 117292
rect 26476 117280 26482 117292
rect 27157 117283 27215 117289
rect 27157 117280 27169 117283
rect 26476 117252 27169 117280
rect 26476 117240 26482 117252
rect 27157 117249 27169 117252
rect 27203 117249 27215 117283
rect 27157 117243 27215 117249
rect 28258 117240 28264 117292
rect 28316 117280 28322 117292
rect 30377 117283 30435 117289
rect 30377 117280 30389 117283
rect 28316 117252 30389 117280
rect 28316 117240 28322 117252
rect 30377 117249 30389 117252
rect 30423 117249 30435 117283
rect 34698 117280 34704 117292
rect 34659 117252 34704 117280
rect 30377 117243 30435 117249
rect 34698 117240 34704 117252
rect 34756 117280 34762 117292
rect 35253 117283 35311 117289
rect 35253 117280 35265 117283
rect 34756 117252 35265 117280
rect 34756 117240 34762 117252
rect 35253 117249 35265 117252
rect 35299 117249 35311 117283
rect 35253 117243 35311 117249
rect 36354 117240 36360 117292
rect 36412 117280 36418 117292
rect 37461 117283 37519 117289
rect 37461 117280 37473 117283
rect 36412 117252 37473 117280
rect 36412 117240 36418 117252
rect 37461 117249 37473 117252
rect 37507 117249 37519 117283
rect 37461 117243 37519 117249
rect 40678 117240 40684 117292
rect 40736 117280 40742 117292
rect 41325 117283 41383 117289
rect 41325 117280 41337 117283
rect 40736 117252 41337 117280
rect 40736 117240 40742 117252
rect 41325 117249 41337 117252
rect 41371 117249 41383 117283
rect 45186 117280 45192 117292
rect 45147 117252 45192 117280
rect 41325 117243 41383 117249
rect 45186 117240 45192 117252
rect 45244 117240 45250 117292
rect 49234 117280 49240 117292
rect 49195 117252 49240 117280
rect 49234 117240 49240 117252
rect 49292 117240 49298 117292
rect 52733 117283 52791 117289
rect 52733 117249 52745 117283
rect 52779 117280 52791 117283
rect 56134 117280 56140 117292
rect 52779 117252 55214 117280
rect 56095 117252 56140 117280
rect 52779 117249 52791 117252
rect 52733 117243 52791 117249
rect 5445 117215 5503 117221
rect 5445 117181 5457 117215
rect 5491 117212 5503 117215
rect 11882 117212 11888 117224
rect 5491 117184 6914 117212
rect 11843 117184 11888 117212
rect 5491 117181 5503 117184
rect 5445 117175 5503 117181
rect 6886 117144 6914 117184
rect 11882 117172 11888 117184
rect 11940 117172 11946 117224
rect 35802 117212 35808 117224
rect 16546 117184 35808 117212
rect 16546 117144 16574 117184
rect 35802 117172 35808 117184
rect 35860 117172 35866 117224
rect 6886 117116 16574 117144
rect 19334 117104 19340 117156
rect 19392 117144 19398 117156
rect 19613 117147 19671 117153
rect 19613 117144 19625 117147
rect 19392 117116 19625 117144
rect 19392 117104 19398 117116
rect 19613 117113 19625 117116
rect 19659 117113 19671 117147
rect 22830 117144 22836 117156
rect 22791 117116 22836 117144
rect 19613 117107 19671 117113
rect 22830 117104 22836 117116
rect 22888 117104 22894 117156
rect 30374 117104 30380 117156
rect 30432 117144 30438 117156
rect 30561 117147 30619 117153
rect 30561 117144 30573 117147
rect 30432 117116 30573 117144
rect 30432 117104 30438 117116
rect 30561 117113 30573 117116
rect 30607 117113 30619 117147
rect 30561 117107 30619 117113
rect 34514 117104 34520 117156
rect 34572 117144 34578 117156
rect 34885 117147 34943 117153
rect 34885 117144 34897 117147
rect 34572 117116 34897 117144
rect 34572 117104 34578 117116
rect 34885 117113 34897 117116
rect 34931 117113 34943 117147
rect 37458 117144 37464 117156
rect 34885 117107 34943 117113
rect 34992 117116 37464 117144
rect 2133 117079 2191 117085
rect 2133 117045 2145 117079
rect 2179 117076 2191 117079
rect 2314 117076 2320 117088
rect 2179 117048 2320 117076
rect 2179 117045 2191 117048
rect 2133 117039 2191 117045
rect 2314 117036 2320 117048
rect 2372 117036 2378 117088
rect 8018 117076 8024 117088
rect 7979 117048 8024 117076
rect 8018 117036 8024 117048
rect 8076 117036 8082 117088
rect 15746 117076 15752 117088
rect 15707 117048 15752 117076
rect 15746 117036 15752 117048
rect 15804 117036 15810 117088
rect 26973 117079 27031 117085
rect 26973 117045 26985 117079
rect 27019 117076 27031 117079
rect 34992 117076 35020 117116
rect 37458 117104 37464 117116
rect 37516 117104 37522 117156
rect 37642 117144 37648 117156
rect 37603 117116 37648 117144
rect 37642 117104 37648 117116
rect 37700 117104 37706 117156
rect 45370 117144 45376 117156
rect 45331 117116 45376 117144
rect 45370 117104 45376 117116
rect 45428 117104 45434 117156
rect 52454 117104 52460 117156
rect 52512 117144 52518 117156
rect 52917 117147 52975 117153
rect 52917 117144 52929 117147
rect 52512 117116 52929 117144
rect 52512 117104 52518 117116
rect 52917 117113 52929 117116
rect 52963 117113 52975 117147
rect 55186 117144 55214 117252
rect 56134 117240 56140 117252
rect 56192 117240 56198 117292
rect 59906 117240 59912 117292
rect 59964 117280 59970 117292
rect 60645 117283 60703 117289
rect 60645 117280 60657 117283
rect 59964 117252 60657 117280
rect 59964 117240 59970 117252
rect 60645 117249 60657 117252
rect 60691 117249 60703 117283
rect 63862 117280 63868 117292
rect 63823 117252 63868 117280
rect 60645 117243 60703 117249
rect 63862 117240 63868 117252
rect 63920 117240 63926 117292
rect 67085 117283 67143 117289
rect 67085 117280 67097 117283
rect 66732 117252 67097 117280
rect 56318 117212 56324 117224
rect 56279 117184 56324 117212
rect 56318 117172 56324 117184
rect 56376 117172 56382 117224
rect 58618 117144 58624 117156
rect 55186 117116 58624 117144
rect 52917 117107 52975 117113
rect 58618 117104 58624 117116
rect 58676 117104 58682 117156
rect 60461 117147 60519 117153
rect 60461 117113 60473 117147
rect 60507 117144 60519 117147
rect 66530 117144 66536 117156
rect 60507 117116 66536 117144
rect 60507 117113 60519 117116
rect 60461 117107 60519 117113
rect 66530 117104 66536 117116
rect 66588 117104 66594 117156
rect 66732 117088 66760 117252
rect 67085 117249 67097 117252
rect 67131 117249 67143 117283
rect 67085 117243 67143 117249
rect 70854 117240 70860 117292
rect 70912 117280 70918 117292
rect 71225 117283 71283 117289
rect 71225 117280 71237 117283
rect 70912 117252 71237 117280
rect 70912 117240 70918 117252
rect 71225 117249 71237 117252
rect 71271 117249 71283 117283
rect 74813 117283 74871 117289
rect 74813 117280 74825 117283
rect 71225 117243 71283 117249
rect 74552 117252 74825 117280
rect 67266 117144 67272 117156
rect 67227 117116 67272 117144
rect 67266 117104 67272 117116
rect 67324 117104 67330 117156
rect 74552 117088 74580 117252
rect 74813 117249 74825 117252
rect 74859 117249 74871 117283
rect 74813 117243 74871 117249
rect 77113 117283 77171 117289
rect 77113 117249 77125 117283
rect 77159 117280 77171 117283
rect 78582 117280 78588 117292
rect 77159 117252 78588 117280
rect 77159 117249 77171 117252
rect 77113 117243 77171 117249
rect 78582 117240 78588 117252
rect 78640 117240 78646 117292
rect 77389 117215 77447 117221
rect 77389 117181 77401 117215
rect 77435 117212 77447 117215
rect 77938 117212 77944 117224
rect 77435 117184 77944 117212
rect 77435 117181 77447 117184
rect 77389 117175 77447 117181
rect 77938 117172 77944 117184
rect 77996 117172 78002 117224
rect 74994 117144 75000 117156
rect 74955 117116 75000 117144
rect 74994 117104 75000 117116
rect 75052 117104 75058 117156
rect 27019 117048 35020 117076
rect 27019 117045 27031 117048
rect 26973 117039 27031 117045
rect 41414 117036 41420 117088
rect 41472 117076 41478 117088
rect 41509 117079 41567 117085
rect 41509 117076 41521 117079
rect 41472 117048 41521 117076
rect 41472 117036 41478 117048
rect 41509 117045 41521 117048
rect 41555 117045 41567 117079
rect 49050 117076 49056 117088
rect 49011 117048 49056 117076
rect 41509 117039 41567 117045
rect 49050 117036 49056 117048
rect 49108 117036 49114 117088
rect 64046 117076 64052 117088
rect 64007 117048 64052 117076
rect 64046 117036 64052 117048
rect 64104 117036 64110 117088
rect 66714 117076 66720 117088
rect 66675 117048 66720 117076
rect 66714 117036 66720 117048
rect 66772 117036 66778 117088
rect 71314 117076 71320 117088
rect 71275 117048 71320 117076
rect 71314 117036 71320 117048
rect 71372 117036 71378 117088
rect 74534 117036 74540 117088
rect 74592 117076 74598 117088
rect 74592 117048 74637 117076
rect 74592 117036 74598 117048
rect 1104 116986 78844 117008
rect 1104 116934 4214 116986
rect 4266 116934 4278 116986
rect 4330 116934 4342 116986
rect 4394 116934 4406 116986
rect 4458 116934 4470 116986
rect 4522 116934 34934 116986
rect 34986 116934 34998 116986
rect 35050 116934 35062 116986
rect 35114 116934 35126 116986
rect 35178 116934 35190 116986
rect 35242 116934 65654 116986
rect 65706 116934 65718 116986
rect 65770 116934 65782 116986
rect 65834 116934 65846 116986
rect 65898 116934 65910 116986
rect 65962 116934 78844 116986
rect 1104 116912 78844 116934
rect 15562 116832 15568 116884
rect 15620 116872 15626 116884
rect 40770 116872 40776 116884
rect 15620 116844 40776 116872
rect 15620 116832 15626 116844
rect 40770 116832 40776 116844
rect 40828 116832 40834 116884
rect 41414 116832 41420 116884
rect 41472 116872 41478 116884
rect 66714 116872 66720 116884
rect 41472 116844 66720 116872
rect 41472 116832 41478 116844
rect 66714 116832 66720 116844
rect 66772 116832 66778 116884
rect 77202 116832 77208 116884
rect 77260 116872 77266 116884
rect 78033 116875 78091 116881
rect 78033 116872 78045 116875
rect 77260 116844 78045 116872
rect 77260 116832 77266 116844
rect 78033 116841 78045 116844
rect 78079 116841 78091 116875
rect 78033 116835 78091 116841
rect 10686 116764 10692 116816
rect 10744 116804 10750 116816
rect 34698 116804 34704 116816
rect 10744 116776 34704 116804
rect 10744 116764 10750 116776
rect 34698 116764 34704 116776
rect 34756 116764 34762 116816
rect 40034 116696 40040 116748
rect 40092 116736 40098 116748
rect 74534 116736 74540 116748
rect 40092 116708 74540 116736
rect 40092 116696 40098 116708
rect 74534 116696 74540 116708
rect 74592 116696 74598 116748
rect 1854 116668 1860 116680
rect 1815 116640 1860 116668
rect 1854 116628 1860 116640
rect 1912 116628 1918 116680
rect 77846 116668 77852 116680
rect 77807 116640 77852 116668
rect 77846 116628 77852 116640
rect 77904 116628 77910 116680
rect 2222 116600 2228 116612
rect 2183 116572 2228 116600
rect 2222 116560 2228 116572
rect 2280 116560 2286 116612
rect 1104 116442 78844 116464
rect 1104 116390 19574 116442
rect 19626 116390 19638 116442
rect 19690 116390 19702 116442
rect 19754 116390 19766 116442
rect 19818 116390 19830 116442
rect 19882 116390 50294 116442
rect 50346 116390 50358 116442
rect 50410 116390 50422 116442
rect 50474 116390 50486 116442
rect 50538 116390 50550 116442
rect 50602 116390 78844 116442
rect 1104 116368 78844 116390
rect 40770 116328 40776 116340
rect 40731 116300 40776 116328
rect 40770 116288 40776 116300
rect 40828 116288 40834 116340
rect 37458 116152 37464 116204
rect 37516 116192 37522 116204
rect 39853 116195 39911 116201
rect 39853 116192 39865 116195
rect 37516 116164 39865 116192
rect 37516 116152 37522 116164
rect 39853 116161 39865 116164
rect 39899 116161 39911 116195
rect 39853 116155 39911 116161
rect 40681 116195 40739 116201
rect 40681 116161 40693 116195
rect 40727 116192 40739 116195
rect 49050 116192 49056 116204
rect 40727 116164 49056 116192
rect 40727 116161 40739 116164
rect 40681 116155 40739 116161
rect 49050 116152 49056 116164
rect 49108 116152 49114 116204
rect 40037 116059 40095 116065
rect 40037 116025 40049 116059
rect 40083 116056 40095 116059
rect 40083 116028 45554 116056
rect 40083 116025 40095 116028
rect 40037 116019 40095 116025
rect 45526 115988 45554 116028
rect 77846 115988 77852 116000
rect 45526 115960 77852 115988
rect 77846 115948 77852 115960
rect 77904 115948 77910 116000
rect 1104 115898 78844 115920
rect 1104 115846 4214 115898
rect 4266 115846 4278 115898
rect 4330 115846 4342 115898
rect 4394 115846 4406 115898
rect 4458 115846 4470 115898
rect 4522 115846 34934 115898
rect 34986 115846 34998 115898
rect 35050 115846 35062 115898
rect 35114 115846 35126 115898
rect 35178 115846 35190 115898
rect 35242 115846 65654 115898
rect 65706 115846 65718 115898
rect 65770 115846 65782 115898
rect 65834 115846 65846 115898
rect 65898 115846 65910 115898
rect 65962 115846 78844 115898
rect 1104 115824 78844 115846
rect 1104 115354 78844 115376
rect 1104 115302 19574 115354
rect 19626 115302 19638 115354
rect 19690 115302 19702 115354
rect 19754 115302 19766 115354
rect 19818 115302 19830 115354
rect 19882 115302 50294 115354
rect 50346 115302 50358 115354
rect 50410 115302 50422 115354
rect 50474 115302 50486 115354
rect 50538 115302 50550 115354
rect 50602 115302 78844 115354
rect 1104 115280 78844 115302
rect 1104 114810 78844 114832
rect 1104 114758 4214 114810
rect 4266 114758 4278 114810
rect 4330 114758 4342 114810
rect 4394 114758 4406 114810
rect 4458 114758 4470 114810
rect 4522 114758 34934 114810
rect 34986 114758 34998 114810
rect 35050 114758 35062 114810
rect 35114 114758 35126 114810
rect 35178 114758 35190 114810
rect 35242 114758 65654 114810
rect 65706 114758 65718 114810
rect 65770 114758 65782 114810
rect 65834 114758 65846 114810
rect 65898 114758 65910 114810
rect 65962 114758 78844 114810
rect 1104 114736 78844 114758
rect 77386 114452 77392 114504
rect 77444 114492 77450 114504
rect 77849 114495 77907 114501
rect 77849 114492 77861 114495
rect 77444 114464 77861 114492
rect 77444 114452 77450 114464
rect 77849 114461 77861 114464
rect 77895 114461 77907 114495
rect 77849 114455 77907 114461
rect 78030 114356 78036 114368
rect 77991 114328 78036 114356
rect 78030 114316 78036 114328
rect 78088 114316 78094 114368
rect 1104 114266 78844 114288
rect 1104 114214 19574 114266
rect 19626 114214 19638 114266
rect 19690 114214 19702 114266
rect 19754 114214 19766 114266
rect 19818 114214 19830 114266
rect 19882 114214 50294 114266
rect 50346 114214 50358 114266
rect 50410 114214 50422 114266
rect 50474 114214 50486 114266
rect 50538 114214 50550 114266
rect 50602 114214 78844 114266
rect 1104 114192 78844 114214
rect 24213 114155 24271 114161
rect 24213 114121 24225 114155
rect 24259 114152 24271 114155
rect 28258 114152 28264 114164
rect 24259 114124 28264 114152
rect 24259 114121 24271 114124
rect 24213 114115 24271 114121
rect 28258 114112 28264 114124
rect 28316 114112 28322 114164
rect 20622 113976 20628 114028
rect 20680 114016 20686 114028
rect 24397 114019 24455 114025
rect 24397 114016 24409 114019
rect 20680 113988 24409 114016
rect 20680 113976 20686 113988
rect 24397 113985 24409 113988
rect 24443 113985 24455 114019
rect 24397 113979 24455 113985
rect 1104 113722 78844 113744
rect 1104 113670 4214 113722
rect 4266 113670 4278 113722
rect 4330 113670 4342 113722
rect 4394 113670 4406 113722
rect 4458 113670 4470 113722
rect 4522 113670 34934 113722
rect 34986 113670 34998 113722
rect 35050 113670 35062 113722
rect 35114 113670 35126 113722
rect 35178 113670 35190 113722
rect 35242 113670 65654 113722
rect 65706 113670 65718 113722
rect 65770 113670 65782 113722
rect 65834 113670 65846 113722
rect 65898 113670 65910 113722
rect 65962 113670 78844 113722
rect 1104 113648 78844 113670
rect 1394 113404 1400 113416
rect 1355 113376 1400 113404
rect 1394 113364 1400 113376
rect 1452 113364 1458 113416
rect 1578 113268 1584 113280
rect 1539 113240 1584 113268
rect 1578 113228 1584 113240
rect 1636 113228 1642 113280
rect 1104 113178 78844 113200
rect 1104 113126 19574 113178
rect 19626 113126 19638 113178
rect 19690 113126 19702 113178
rect 19754 113126 19766 113178
rect 19818 113126 19830 113178
rect 19882 113126 50294 113178
rect 50346 113126 50358 113178
rect 50410 113126 50422 113178
rect 50474 113126 50486 113178
rect 50538 113126 50550 113178
rect 50602 113126 78844 113178
rect 1104 113104 78844 113126
rect 1104 112634 78844 112656
rect 1104 112582 4214 112634
rect 4266 112582 4278 112634
rect 4330 112582 4342 112634
rect 4394 112582 4406 112634
rect 4458 112582 4470 112634
rect 4522 112582 34934 112634
rect 34986 112582 34998 112634
rect 35050 112582 35062 112634
rect 35114 112582 35126 112634
rect 35178 112582 35190 112634
rect 35242 112582 65654 112634
rect 65706 112582 65718 112634
rect 65770 112582 65782 112634
rect 65834 112582 65846 112634
rect 65898 112582 65910 112634
rect 65962 112582 78844 112634
rect 1104 112560 78844 112582
rect 1104 112090 78844 112112
rect 1104 112038 19574 112090
rect 19626 112038 19638 112090
rect 19690 112038 19702 112090
rect 19754 112038 19766 112090
rect 19818 112038 19830 112090
rect 19882 112038 50294 112090
rect 50346 112038 50358 112090
rect 50410 112038 50422 112090
rect 50474 112038 50486 112090
rect 50538 112038 50550 112090
rect 50602 112038 78844 112090
rect 1104 112016 78844 112038
rect 66530 111908 66536 111920
rect 66491 111880 66536 111908
rect 66530 111868 66536 111880
rect 66588 111868 66594 111920
rect 66717 111843 66775 111849
rect 66717 111809 66729 111843
rect 66763 111840 66775 111843
rect 76006 111840 76012 111852
rect 66763 111812 76012 111840
rect 66763 111809 66775 111812
rect 66717 111803 66775 111809
rect 76006 111800 76012 111812
rect 76064 111800 76070 111852
rect 1104 111546 78844 111568
rect 1104 111494 4214 111546
rect 4266 111494 4278 111546
rect 4330 111494 4342 111546
rect 4394 111494 4406 111546
rect 4458 111494 4470 111546
rect 4522 111494 34934 111546
rect 34986 111494 34998 111546
rect 35050 111494 35062 111546
rect 35114 111494 35126 111546
rect 35178 111494 35190 111546
rect 35242 111494 65654 111546
rect 65706 111494 65718 111546
rect 65770 111494 65782 111546
rect 65834 111494 65846 111546
rect 65898 111494 65910 111546
rect 65962 111494 78844 111546
rect 1104 111472 78844 111494
rect 1104 111002 78844 111024
rect 1104 110950 19574 111002
rect 19626 110950 19638 111002
rect 19690 110950 19702 111002
rect 19754 110950 19766 111002
rect 19818 110950 19830 111002
rect 19882 110950 50294 111002
rect 50346 110950 50358 111002
rect 50410 110950 50422 111002
rect 50474 110950 50486 111002
rect 50538 110950 50550 111002
rect 50602 110950 78844 111002
rect 1104 110928 78844 110950
rect 77665 110755 77723 110761
rect 77665 110721 77677 110755
rect 77711 110752 77723 110755
rect 77754 110752 77760 110764
rect 77711 110724 77760 110752
rect 77711 110721 77723 110724
rect 77665 110715 77723 110721
rect 77754 110712 77760 110724
rect 77812 110712 77818 110764
rect 77846 110548 77852 110560
rect 77807 110520 77852 110548
rect 77846 110508 77852 110520
rect 77904 110508 77910 110560
rect 1104 110458 78844 110480
rect 1104 110406 4214 110458
rect 4266 110406 4278 110458
rect 4330 110406 4342 110458
rect 4394 110406 4406 110458
rect 4458 110406 4470 110458
rect 4522 110406 34934 110458
rect 34986 110406 34998 110458
rect 35050 110406 35062 110458
rect 35114 110406 35126 110458
rect 35178 110406 35190 110458
rect 35242 110406 65654 110458
rect 65706 110406 65718 110458
rect 65770 110406 65782 110458
rect 65834 110406 65846 110458
rect 65898 110406 65910 110458
rect 65962 110406 78844 110458
rect 1104 110384 78844 110406
rect 1104 109914 78844 109936
rect 1104 109862 19574 109914
rect 19626 109862 19638 109914
rect 19690 109862 19702 109914
rect 19754 109862 19766 109914
rect 19818 109862 19830 109914
rect 19882 109862 50294 109914
rect 50346 109862 50358 109914
rect 50410 109862 50422 109914
rect 50474 109862 50486 109914
rect 50538 109862 50550 109914
rect 50602 109862 78844 109914
rect 1104 109840 78844 109862
rect 1854 109664 1860 109676
rect 1815 109636 1860 109664
rect 1854 109624 1860 109636
rect 1912 109624 1918 109676
rect 1949 109463 2007 109469
rect 1949 109429 1961 109463
rect 1995 109460 2007 109463
rect 20622 109460 20628 109472
rect 1995 109432 20628 109460
rect 1995 109429 2007 109432
rect 1949 109423 2007 109429
rect 20622 109420 20628 109432
rect 20680 109420 20686 109472
rect 1104 109370 78844 109392
rect 1104 109318 4214 109370
rect 4266 109318 4278 109370
rect 4330 109318 4342 109370
rect 4394 109318 4406 109370
rect 4458 109318 4470 109370
rect 4522 109318 34934 109370
rect 34986 109318 34998 109370
rect 35050 109318 35062 109370
rect 35114 109318 35126 109370
rect 35178 109318 35190 109370
rect 35242 109318 65654 109370
rect 65706 109318 65718 109370
rect 65770 109318 65782 109370
rect 65834 109318 65846 109370
rect 65898 109318 65910 109370
rect 65962 109318 78844 109370
rect 1104 109296 78844 109318
rect 40034 109256 40040 109268
rect 39995 109228 40040 109256
rect 40034 109216 40040 109228
rect 40092 109216 40098 109268
rect 39850 109052 39856 109064
rect 39811 109024 39856 109052
rect 39850 109012 39856 109024
rect 39908 109012 39914 109064
rect 1104 108826 78844 108848
rect 1104 108774 19574 108826
rect 19626 108774 19638 108826
rect 19690 108774 19702 108826
rect 19754 108774 19766 108826
rect 19818 108774 19830 108826
rect 19882 108774 50294 108826
rect 50346 108774 50358 108826
rect 50410 108774 50422 108826
rect 50474 108774 50486 108826
rect 50538 108774 50550 108826
rect 50602 108774 78844 108826
rect 1104 108752 78844 108774
rect 1104 108282 78844 108304
rect 1104 108230 4214 108282
rect 4266 108230 4278 108282
rect 4330 108230 4342 108282
rect 4394 108230 4406 108282
rect 4458 108230 4470 108282
rect 4522 108230 34934 108282
rect 34986 108230 34998 108282
rect 35050 108230 35062 108282
rect 35114 108230 35126 108282
rect 35178 108230 35190 108282
rect 35242 108230 65654 108282
rect 65706 108230 65718 108282
rect 65770 108230 65782 108282
rect 65834 108230 65846 108282
rect 65898 108230 65910 108282
rect 65962 108230 78844 108282
rect 1104 108208 78844 108230
rect 1104 107738 78844 107760
rect 1104 107686 19574 107738
rect 19626 107686 19638 107738
rect 19690 107686 19702 107738
rect 19754 107686 19766 107738
rect 19818 107686 19830 107738
rect 19882 107686 50294 107738
rect 50346 107686 50358 107738
rect 50410 107686 50422 107738
rect 50474 107686 50486 107738
rect 50538 107686 50550 107738
rect 50602 107686 78844 107738
rect 1104 107664 78844 107686
rect 1104 107194 78844 107216
rect 1104 107142 4214 107194
rect 4266 107142 4278 107194
rect 4330 107142 4342 107194
rect 4394 107142 4406 107194
rect 4458 107142 4470 107194
rect 4522 107142 34934 107194
rect 34986 107142 34998 107194
rect 35050 107142 35062 107194
rect 35114 107142 35126 107194
rect 35178 107142 35190 107194
rect 35242 107142 65654 107194
rect 65706 107142 65718 107194
rect 65770 107142 65782 107194
rect 65834 107142 65846 107194
rect 65898 107142 65910 107194
rect 65962 107142 78844 107194
rect 1104 107120 78844 107142
rect 1104 106650 78844 106672
rect 1104 106598 19574 106650
rect 19626 106598 19638 106650
rect 19690 106598 19702 106650
rect 19754 106598 19766 106650
rect 19818 106598 19830 106650
rect 19882 106598 50294 106650
rect 50346 106598 50358 106650
rect 50410 106598 50422 106650
rect 50474 106598 50486 106650
rect 50538 106598 50550 106650
rect 50602 106598 78844 106650
rect 1104 106576 78844 106598
rect 76006 106360 76012 106412
rect 76064 106400 76070 106412
rect 77665 106403 77723 106409
rect 77665 106400 77677 106403
rect 76064 106372 77677 106400
rect 76064 106360 76070 106372
rect 77665 106369 77677 106372
rect 77711 106369 77723 106403
rect 77665 106363 77723 106369
rect 77846 106196 77852 106208
rect 77807 106168 77852 106196
rect 77846 106156 77852 106168
rect 77904 106156 77910 106208
rect 1104 106106 78844 106128
rect 1104 106054 4214 106106
rect 4266 106054 4278 106106
rect 4330 106054 4342 106106
rect 4394 106054 4406 106106
rect 4458 106054 4470 106106
rect 4522 106054 34934 106106
rect 34986 106054 34998 106106
rect 35050 106054 35062 106106
rect 35114 106054 35126 106106
rect 35178 106054 35190 106106
rect 35242 106054 65654 106106
rect 65706 106054 65718 106106
rect 65770 106054 65782 106106
rect 65834 106054 65846 106106
rect 65898 106054 65910 106106
rect 65962 106054 78844 106106
rect 1104 106032 78844 106054
rect 1394 105788 1400 105800
rect 1355 105760 1400 105788
rect 1394 105748 1400 105760
rect 1452 105748 1458 105800
rect 1673 105723 1731 105729
rect 1673 105689 1685 105723
rect 1719 105720 1731 105723
rect 1854 105720 1860 105732
rect 1719 105692 1860 105720
rect 1719 105689 1731 105692
rect 1673 105683 1731 105689
rect 1854 105680 1860 105692
rect 1912 105680 1918 105732
rect 1104 105562 78844 105584
rect 1104 105510 19574 105562
rect 19626 105510 19638 105562
rect 19690 105510 19702 105562
rect 19754 105510 19766 105562
rect 19818 105510 19830 105562
rect 19882 105510 50294 105562
rect 50346 105510 50358 105562
rect 50410 105510 50422 105562
rect 50474 105510 50486 105562
rect 50538 105510 50550 105562
rect 50602 105510 78844 105562
rect 1104 105488 78844 105510
rect 1104 105018 78844 105040
rect 1104 104966 4214 105018
rect 4266 104966 4278 105018
rect 4330 104966 4342 105018
rect 4394 104966 4406 105018
rect 4458 104966 4470 105018
rect 4522 104966 34934 105018
rect 34986 104966 34998 105018
rect 35050 104966 35062 105018
rect 35114 104966 35126 105018
rect 35178 104966 35190 105018
rect 35242 104966 65654 105018
rect 65706 104966 65718 105018
rect 65770 104966 65782 105018
rect 65834 104966 65846 105018
rect 65898 104966 65910 105018
rect 65962 104966 78844 105018
rect 1104 104944 78844 104966
rect 1104 104474 78844 104496
rect 1104 104422 19574 104474
rect 19626 104422 19638 104474
rect 19690 104422 19702 104474
rect 19754 104422 19766 104474
rect 19818 104422 19830 104474
rect 19882 104422 50294 104474
rect 50346 104422 50358 104474
rect 50410 104422 50422 104474
rect 50474 104422 50486 104474
rect 50538 104422 50550 104474
rect 50602 104422 78844 104474
rect 1104 104400 78844 104422
rect 1104 103930 78844 103952
rect 1104 103878 4214 103930
rect 4266 103878 4278 103930
rect 4330 103878 4342 103930
rect 4394 103878 4406 103930
rect 4458 103878 4470 103930
rect 4522 103878 34934 103930
rect 34986 103878 34998 103930
rect 35050 103878 35062 103930
rect 35114 103878 35126 103930
rect 35178 103878 35190 103930
rect 35242 103878 65654 103930
rect 65706 103878 65718 103930
rect 65770 103878 65782 103930
rect 65834 103878 65846 103930
rect 65898 103878 65910 103930
rect 65962 103878 78844 103930
rect 1104 103856 78844 103878
rect 77849 103751 77907 103757
rect 77849 103717 77861 103751
rect 77895 103748 77907 103751
rect 77938 103748 77944 103760
rect 77895 103720 77944 103748
rect 77895 103717 77907 103720
rect 77849 103711 77907 103717
rect 77938 103708 77944 103720
rect 77996 103708 78002 103760
rect 78030 103612 78036 103624
rect 77991 103584 78036 103612
rect 78030 103572 78036 103584
rect 78088 103572 78094 103624
rect 1104 103386 78844 103408
rect 1104 103334 19574 103386
rect 19626 103334 19638 103386
rect 19690 103334 19702 103386
rect 19754 103334 19766 103386
rect 19818 103334 19830 103386
rect 19882 103334 50294 103386
rect 50346 103334 50358 103386
rect 50410 103334 50422 103386
rect 50474 103334 50486 103386
rect 50538 103334 50550 103386
rect 50602 103334 78844 103386
rect 1104 103312 78844 103334
rect 77294 103096 77300 103148
rect 77352 103136 77358 103148
rect 77665 103139 77723 103145
rect 77665 103136 77677 103139
rect 77352 103108 77677 103136
rect 77352 103096 77358 103108
rect 77665 103105 77677 103108
rect 77711 103105 77723 103139
rect 77665 103099 77723 103105
rect 77294 102932 77300 102944
rect 77255 102904 77300 102932
rect 77294 102892 77300 102904
rect 77352 102892 77358 102944
rect 77846 102932 77852 102944
rect 77807 102904 77852 102932
rect 77846 102892 77852 102904
rect 77904 102892 77910 102944
rect 1104 102842 78844 102864
rect 1104 102790 4214 102842
rect 4266 102790 4278 102842
rect 4330 102790 4342 102842
rect 4394 102790 4406 102842
rect 4458 102790 4470 102842
rect 4522 102790 34934 102842
rect 34986 102790 34998 102842
rect 35050 102790 35062 102842
rect 35114 102790 35126 102842
rect 35178 102790 35190 102842
rect 35242 102790 65654 102842
rect 65706 102790 65718 102842
rect 65770 102790 65782 102842
rect 65834 102790 65846 102842
rect 65898 102790 65910 102842
rect 65962 102790 78844 102842
rect 1104 102768 78844 102790
rect 1104 102298 78844 102320
rect 1104 102246 19574 102298
rect 19626 102246 19638 102298
rect 19690 102246 19702 102298
rect 19754 102246 19766 102298
rect 19818 102246 19830 102298
rect 19882 102246 50294 102298
rect 50346 102246 50358 102298
rect 50410 102246 50422 102298
rect 50474 102246 50486 102298
rect 50538 102246 50550 102298
rect 50602 102246 78844 102298
rect 1104 102224 78844 102246
rect 1104 101754 78844 101776
rect 1104 101702 4214 101754
rect 4266 101702 4278 101754
rect 4330 101702 4342 101754
rect 4394 101702 4406 101754
rect 4458 101702 4470 101754
rect 4522 101702 34934 101754
rect 34986 101702 34998 101754
rect 35050 101702 35062 101754
rect 35114 101702 35126 101754
rect 35178 101702 35190 101754
rect 35242 101702 65654 101754
rect 65706 101702 65718 101754
rect 65770 101702 65782 101754
rect 65834 101702 65846 101754
rect 65898 101702 65910 101754
rect 65962 101702 78844 101754
rect 1104 101680 78844 101702
rect 1394 101436 1400 101448
rect 1355 101408 1400 101436
rect 1394 101396 1400 101408
rect 1452 101396 1458 101448
rect 1581 101303 1639 101309
rect 1581 101269 1593 101303
rect 1627 101300 1639 101303
rect 39850 101300 39856 101312
rect 1627 101272 39856 101300
rect 1627 101269 1639 101272
rect 1581 101263 1639 101269
rect 39850 101260 39856 101272
rect 39908 101260 39914 101312
rect 1104 101210 78844 101232
rect 1104 101158 19574 101210
rect 19626 101158 19638 101210
rect 19690 101158 19702 101210
rect 19754 101158 19766 101210
rect 19818 101158 19830 101210
rect 19882 101158 50294 101210
rect 50346 101158 50358 101210
rect 50410 101158 50422 101210
rect 50474 101158 50486 101210
rect 50538 101158 50550 101210
rect 50602 101158 78844 101210
rect 1104 101136 78844 101158
rect 1104 100666 78844 100688
rect 1104 100614 4214 100666
rect 4266 100614 4278 100666
rect 4330 100614 4342 100666
rect 4394 100614 4406 100666
rect 4458 100614 4470 100666
rect 4522 100614 34934 100666
rect 34986 100614 34998 100666
rect 35050 100614 35062 100666
rect 35114 100614 35126 100666
rect 35178 100614 35190 100666
rect 35242 100614 65654 100666
rect 65706 100614 65718 100666
rect 65770 100614 65782 100666
rect 65834 100614 65846 100666
rect 65898 100614 65910 100666
rect 65962 100614 78844 100666
rect 1104 100592 78844 100614
rect 58618 100552 58624 100564
rect 58579 100524 58624 100552
rect 58618 100512 58624 100524
rect 58676 100512 58682 100564
rect 58526 100280 58532 100292
rect 58487 100252 58532 100280
rect 58526 100240 58532 100252
rect 58584 100240 58590 100292
rect 1104 100122 78844 100144
rect 1104 100070 19574 100122
rect 19626 100070 19638 100122
rect 19690 100070 19702 100122
rect 19754 100070 19766 100122
rect 19818 100070 19830 100122
rect 19882 100070 50294 100122
rect 50346 100070 50358 100122
rect 50410 100070 50422 100122
rect 50474 100070 50486 100122
rect 50538 100070 50550 100122
rect 50602 100070 78844 100122
rect 1104 100048 78844 100070
rect 1104 99578 78844 99600
rect 1104 99526 4214 99578
rect 4266 99526 4278 99578
rect 4330 99526 4342 99578
rect 4394 99526 4406 99578
rect 4458 99526 4470 99578
rect 4522 99526 34934 99578
rect 34986 99526 34998 99578
rect 35050 99526 35062 99578
rect 35114 99526 35126 99578
rect 35178 99526 35190 99578
rect 35242 99526 65654 99578
rect 65706 99526 65718 99578
rect 65770 99526 65782 99578
rect 65834 99526 65846 99578
rect 65898 99526 65910 99578
rect 65962 99526 78844 99578
rect 1104 99504 78844 99526
rect 1104 99034 78844 99056
rect 1104 98982 19574 99034
rect 19626 98982 19638 99034
rect 19690 98982 19702 99034
rect 19754 98982 19766 99034
rect 19818 98982 19830 99034
rect 19882 98982 50294 99034
rect 50346 98982 50358 99034
rect 50410 98982 50422 99034
rect 50474 98982 50486 99034
rect 50538 98982 50550 99034
rect 50602 98982 78844 99034
rect 1104 98960 78844 98982
rect 77665 98787 77723 98793
rect 77665 98753 77677 98787
rect 77711 98784 77723 98787
rect 78122 98784 78128 98796
rect 77711 98756 78128 98784
rect 77711 98753 77723 98756
rect 77665 98747 77723 98753
rect 78122 98744 78128 98756
rect 78180 98744 78186 98796
rect 77846 98648 77852 98660
rect 77807 98620 77852 98648
rect 77846 98608 77852 98620
rect 77904 98608 77910 98660
rect 1104 98490 78844 98512
rect 1104 98438 4214 98490
rect 4266 98438 4278 98490
rect 4330 98438 4342 98490
rect 4394 98438 4406 98490
rect 4458 98438 4470 98490
rect 4522 98438 34934 98490
rect 34986 98438 34998 98490
rect 35050 98438 35062 98490
rect 35114 98438 35126 98490
rect 35178 98438 35190 98490
rect 35242 98438 65654 98490
rect 65706 98438 65718 98490
rect 65770 98438 65782 98490
rect 65834 98438 65846 98490
rect 65898 98438 65910 98490
rect 65962 98438 78844 98490
rect 1104 98416 78844 98438
rect 1104 97946 78844 97968
rect 1104 97894 19574 97946
rect 19626 97894 19638 97946
rect 19690 97894 19702 97946
rect 19754 97894 19766 97946
rect 19818 97894 19830 97946
rect 19882 97894 50294 97946
rect 50346 97894 50358 97946
rect 50410 97894 50422 97946
rect 50474 97894 50486 97946
rect 50538 97894 50550 97946
rect 50602 97894 78844 97946
rect 1104 97872 78844 97894
rect 1394 97696 1400 97708
rect 1355 97668 1400 97696
rect 1394 97656 1400 97668
rect 1452 97656 1458 97708
rect 1670 97628 1676 97640
rect 1631 97600 1676 97628
rect 1670 97588 1676 97600
rect 1728 97588 1734 97640
rect 1104 97402 78844 97424
rect 1104 97350 4214 97402
rect 4266 97350 4278 97402
rect 4330 97350 4342 97402
rect 4394 97350 4406 97402
rect 4458 97350 4470 97402
rect 4522 97350 34934 97402
rect 34986 97350 34998 97402
rect 35050 97350 35062 97402
rect 35114 97350 35126 97402
rect 35178 97350 35190 97402
rect 35242 97350 65654 97402
rect 65706 97350 65718 97402
rect 65770 97350 65782 97402
rect 65834 97350 65846 97402
rect 65898 97350 65910 97402
rect 65962 97350 78844 97402
rect 1104 97328 78844 97350
rect 1104 96858 78844 96880
rect 1104 96806 19574 96858
rect 19626 96806 19638 96858
rect 19690 96806 19702 96858
rect 19754 96806 19766 96858
rect 19818 96806 19830 96858
rect 19882 96806 50294 96858
rect 50346 96806 50358 96858
rect 50410 96806 50422 96858
rect 50474 96806 50486 96858
rect 50538 96806 50550 96858
rect 50602 96806 78844 96858
rect 1104 96784 78844 96806
rect 1104 96314 78844 96336
rect 1104 96262 4214 96314
rect 4266 96262 4278 96314
rect 4330 96262 4342 96314
rect 4394 96262 4406 96314
rect 4458 96262 4470 96314
rect 4522 96262 34934 96314
rect 34986 96262 34998 96314
rect 35050 96262 35062 96314
rect 35114 96262 35126 96314
rect 35178 96262 35190 96314
rect 35242 96262 65654 96314
rect 65706 96262 65718 96314
rect 65770 96262 65782 96314
rect 65834 96262 65846 96314
rect 65898 96262 65910 96314
rect 65962 96262 78844 96314
rect 1104 96240 78844 96262
rect 40310 95928 40316 95940
rect 40271 95900 40316 95928
rect 40310 95888 40316 95900
rect 40368 95888 40374 95940
rect 1486 95820 1492 95872
rect 1544 95860 1550 95872
rect 40405 95863 40463 95869
rect 40405 95860 40417 95863
rect 1544 95832 40417 95860
rect 1544 95820 1550 95832
rect 40405 95829 40417 95832
rect 40451 95829 40463 95863
rect 40405 95823 40463 95829
rect 1104 95770 78844 95792
rect 1104 95718 19574 95770
rect 19626 95718 19638 95770
rect 19690 95718 19702 95770
rect 19754 95718 19766 95770
rect 19818 95718 19830 95770
rect 19882 95718 50294 95770
rect 50346 95718 50358 95770
rect 50410 95718 50422 95770
rect 50474 95718 50486 95770
rect 50538 95718 50550 95770
rect 50602 95718 78844 95770
rect 1104 95696 78844 95718
rect 1104 95226 78844 95248
rect 1104 95174 4214 95226
rect 4266 95174 4278 95226
rect 4330 95174 4342 95226
rect 4394 95174 4406 95226
rect 4458 95174 4470 95226
rect 4522 95174 34934 95226
rect 34986 95174 34998 95226
rect 35050 95174 35062 95226
rect 35114 95174 35126 95226
rect 35178 95174 35190 95226
rect 35242 95174 65654 95226
rect 65706 95174 65718 95226
rect 65770 95174 65782 95226
rect 65834 95174 65846 95226
rect 65898 95174 65910 95226
rect 65962 95174 78844 95226
rect 1104 95152 78844 95174
rect 77849 94911 77907 94917
rect 77849 94877 77861 94911
rect 77895 94908 77907 94911
rect 77938 94908 77944 94920
rect 77895 94880 77944 94908
rect 77895 94877 77907 94880
rect 77849 94871 77907 94877
rect 77938 94868 77944 94880
rect 77996 94868 78002 94920
rect 78030 94772 78036 94784
rect 77991 94744 78036 94772
rect 78030 94732 78036 94744
rect 78088 94732 78094 94784
rect 1104 94682 78844 94704
rect 1104 94630 19574 94682
rect 19626 94630 19638 94682
rect 19690 94630 19702 94682
rect 19754 94630 19766 94682
rect 19818 94630 19830 94682
rect 19882 94630 50294 94682
rect 50346 94630 50358 94682
rect 50410 94630 50422 94682
rect 50474 94630 50486 94682
rect 50538 94630 50550 94682
rect 50602 94630 78844 94682
rect 1104 94608 78844 94630
rect 1397 94435 1455 94441
rect 1397 94401 1409 94435
rect 1443 94432 1455 94435
rect 2958 94432 2964 94444
rect 1443 94404 2964 94432
rect 1443 94401 1455 94404
rect 1397 94395 1455 94401
rect 2958 94392 2964 94404
rect 3016 94392 3022 94444
rect 1578 94228 1584 94240
rect 1539 94200 1584 94228
rect 1578 94188 1584 94200
rect 1636 94188 1642 94240
rect 1104 94138 78844 94160
rect 1104 94086 4214 94138
rect 4266 94086 4278 94138
rect 4330 94086 4342 94138
rect 4394 94086 4406 94138
rect 4458 94086 4470 94138
rect 4522 94086 34934 94138
rect 34986 94086 34998 94138
rect 35050 94086 35062 94138
rect 35114 94086 35126 94138
rect 35178 94086 35190 94138
rect 35242 94086 65654 94138
rect 65706 94086 65718 94138
rect 65770 94086 65782 94138
rect 65834 94086 65846 94138
rect 65898 94086 65910 94138
rect 65962 94086 78844 94138
rect 1104 94064 78844 94086
rect 1104 93594 78844 93616
rect 1104 93542 19574 93594
rect 19626 93542 19638 93594
rect 19690 93542 19702 93594
rect 19754 93542 19766 93594
rect 19818 93542 19830 93594
rect 19882 93542 50294 93594
rect 50346 93542 50358 93594
rect 50410 93542 50422 93594
rect 50474 93542 50486 93594
rect 50538 93542 50550 93594
rect 50602 93542 78844 93594
rect 1104 93520 78844 93542
rect 1104 93050 78844 93072
rect 1104 92998 4214 93050
rect 4266 92998 4278 93050
rect 4330 92998 4342 93050
rect 4394 92998 4406 93050
rect 4458 92998 4470 93050
rect 4522 92998 34934 93050
rect 34986 92998 34998 93050
rect 35050 92998 35062 93050
rect 35114 92998 35126 93050
rect 35178 92998 35190 93050
rect 35242 92998 65654 93050
rect 65706 92998 65718 93050
rect 65770 92998 65782 93050
rect 65834 92998 65846 93050
rect 65898 92998 65910 93050
rect 65962 92998 78844 93050
rect 1104 92976 78844 92998
rect 1104 92506 78844 92528
rect 1104 92454 19574 92506
rect 19626 92454 19638 92506
rect 19690 92454 19702 92506
rect 19754 92454 19766 92506
rect 19818 92454 19830 92506
rect 19882 92454 50294 92506
rect 50346 92454 50358 92506
rect 50410 92454 50422 92506
rect 50474 92454 50486 92506
rect 50538 92454 50550 92506
rect 50602 92454 78844 92506
rect 1104 92432 78844 92454
rect 41414 92392 41420 92404
rect 41375 92364 41420 92392
rect 41414 92352 41420 92364
rect 41472 92352 41478 92404
rect 41046 92216 41052 92268
rect 41104 92256 41110 92268
rect 41325 92259 41383 92265
rect 41325 92256 41337 92259
rect 41104 92228 41337 92256
rect 41104 92216 41110 92228
rect 41325 92225 41337 92228
rect 41371 92225 41383 92259
rect 41325 92219 41383 92225
rect 1104 91962 78844 91984
rect 1104 91910 4214 91962
rect 4266 91910 4278 91962
rect 4330 91910 4342 91962
rect 4394 91910 4406 91962
rect 4458 91910 4470 91962
rect 4522 91910 34934 91962
rect 34986 91910 34998 91962
rect 35050 91910 35062 91962
rect 35114 91910 35126 91962
rect 35178 91910 35190 91962
rect 35242 91910 65654 91962
rect 65706 91910 65718 91962
rect 65770 91910 65782 91962
rect 65834 91910 65846 91962
rect 65898 91910 65910 91962
rect 65962 91910 78844 91962
rect 1104 91888 78844 91910
rect 1104 91418 78844 91440
rect 1104 91366 19574 91418
rect 19626 91366 19638 91418
rect 19690 91366 19702 91418
rect 19754 91366 19766 91418
rect 19818 91366 19830 91418
rect 19882 91366 50294 91418
rect 50346 91366 50358 91418
rect 50410 91366 50422 91418
rect 50474 91366 50486 91418
rect 50538 91366 50550 91418
rect 50602 91366 78844 91418
rect 1104 91344 78844 91366
rect 1104 90874 78844 90896
rect 1104 90822 4214 90874
rect 4266 90822 4278 90874
rect 4330 90822 4342 90874
rect 4394 90822 4406 90874
rect 4458 90822 4470 90874
rect 4522 90822 34934 90874
rect 34986 90822 34998 90874
rect 35050 90822 35062 90874
rect 35114 90822 35126 90874
rect 35178 90822 35190 90874
rect 35242 90822 65654 90874
rect 65706 90822 65718 90874
rect 65770 90822 65782 90874
rect 65834 90822 65846 90874
rect 65898 90822 65910 90874
rect 65962 90822 78844 90874
rect 1104 90800 78844 90822
rect 77938 90488 77944 90500
rect 77899 90460 77944 90488
rect 77938 90448 77944 90460
rect 77996 90448 78002 90500
rect 58526 90380 58532 90432
rect 58584 90420 58590 90432
rect 78033 90423 78091 90429
rect 78033 90420 78045 90423
rect 58584 90392 78045 90420
rect 58584 90380 58590 90392
rect 78033 90389 78045 90392
rect 78079 90389 78091 90423
rect 78033 90383 78091 90389
rect 1104 90330 78844 90352
rect 1104 90278 19574 90330
rect 19626 90278 19638 90330
rect 19690 90278 19702 90330
rect 19754 90278 19766 90330
rect 19818 90278 19830 90330
rect 19882 90278 50294 90330
rect 50346 90278 50358 90330
rect 50410 90278 50422 90330
rect 50474 90278 50486 90330
rect 50538 90278 50550 90330
rect 50602 90278 78844 90330
rect 1104 90256 78844 90278
rect 1486 90080 1492 90092
rect 1447 90052 1492 90080
rect 1486 90040 1492 90052
rect 1544 90040 1550 90092
rect 2041 90015 2099 90021
rect 2041 89981 2053 90015
rect 2087 90012 2099 90015
rect 41046 90012 41052 90024
rect 2087 89984 41052 90012
rect 2087 89981 2099 89984
rect 2041 89975 2099 89981
rect 41046 89972 41052 89984
rect 41104 89972 41110 90024
rect 1104 89786 78844 89808
rect 1104 89734 4214 89786
rect 4266 89734 4278 89786
rect 4330 89734 4342 89786
rect 4394 89734 4406 89786
rect 4458 89734 4470 89786
rect 4522 89734 34934 89786
rect 34986 89734 34998 89786
rect 35050 89734 35062 89786
rect 35114 89734 35126 89786
rect 35178 89734 35190 89786
rect 35242 89734 65654 89786
rect 65706 89734 65718 89786
rect 65770 89734 65782 89786
rect 65834 89734 65846 89786
rect 65898 89734 65910 89786
rect 65962 89734 78844 89786
rect 1104 89712 78844 89734
rect 1104 89242 78844 89264
rect 1104 89190 19574 89242
rect 19626 89190 19638 89242
rect 19690 89190 19702 89242
rect 19754 89190 19766 89242
rect 19818 89190 19830 89242
rect 19882 89190 50294 89242
rect 50346 89190 50358 89242
rect 50410 89190 50422 89242
rect 50474 89190 50486 89242
rect 50538 89190 50550 89242
rect 50602 89190 78844 89242
rect 1104 89168 78844 89190
rect 39942 88992 39948 89004
rect 39903 88964 39948 88992
rect 39942 88952 39948 88964
rect 40000 88952 40006 89004
rect 7834 88748 7840 88800
rect 7892 88788 7898 88800
rect 40037 88791 40095 88797
rect 40037 88788 40049 88791
rect 7892 88760 40049 88788
rect 7892 88748 7898 88760
rect 40037 88757 40049 88760
rect 40083 88757 40095 88791
rect 40037 88751 40095 88757
rect 1104 88698 78844 88720
rect 1104 88646 4214 88698
rect 4266 88646 4278 88698
rect 4330 88646 4342 88698
rect 4394 88646 4406 88698
rect 4458 88646 4470 88698
rect 4522 88646 34934 88698
rect 34986 88646 34998 88698
rect 35050 88646 35062 88698
rect 35114 88646 35126 88698
rect 35178 88646 35190 88698
rect 35242 88646 65654 88698
rect 65706 88646 65718 88698
rect 65770 88646 65782 88698
rect 65834 88646 65846 88698
rect 65898 88646 65910 88698
rect 65962 88646 78844 88698
rect 1104 88624 78844 88646
rect 1104 88154 78844 88176
rect 1104 88102 19574 88154
rect 19626 88102 19638 88154
rect 19690 88102 19702 88154
rect 19754 88102 19766 88154
rect 19818 88102 19830 88154
rect 19882 88102 50294 88154
rect 50346 88102 50358 88154
rect 50410 88102 50422 88154
rect 50474 88102 50486 88154
rect 50538 88102 50550 88154
rect 50602 88102 78844 88154
rect 1104 88080 78844 88102
rect 1104 87610 78844 87632
rect 1104 87558 4214 87610
rect 4266 87558 4278 87610
rect 4330 87558 4342 87610
rect 4394 87558 4406 87610
rect 4458 87558 4470 87610
rect 4522 87558 34934 87610
rect 34986 87558 34998 87610
rect 35050 87558 35062 87610
rect 35114 87558 35126 87610
rect 35178 87558 35190 87610
rect 35242 87558 65654 87610
rect 65706 87558 65718 87610
rect 65770 87558 65782 87610
rect 65834 87558 65846 87610
rect 65898 87558 65910 87610
rect 65962 87558 78844 87610
rect 1104 87536 78844 87558
rect 77757 87227 77815 87233
rect 77757 87193 77769 87227
rect 77803 87224 77815 87227
rect 77938 87224 77944 87236
rect 77803 87196 77944 87224
rect 77803 87193 77815 87196
rect 77757 87187 77815 87193
rect 77938 87184 77944 87196
rect 77996 87184 78002 87236
rect 40310 87116 40316 87168
rect 40368 87156 40374 87168
rect 77849 87159 77907 87165
rect 77849 87156 77861 87159
rect 40368 87128 77861 87156
rect 40368 87116 40374 87128
rect 77849 87125 77861 87128
rect 77895 87125 77907 87159
rect 77849 87119 77907 87125
rect 1104 87066 78844 87088
rect 1104 87014 19574 87066
rect 19626 87014 19638 87066
rect 19690 87014 19702 87066
rect 19754 87014 19766 87066
rect 19818 87014 19830 87066
rect 19882 87014 50294 87066
rect 50346 87014 50358 87066
rect 50410 87014 50422 87066
rect 50474 87014 50486 87066
rect 50538 87014 50550 87066
rect 50602 87014 78844 87066
rect 1104 86992 78844 87014
rect 1104 86522 78844 86544
rect 1104 86470 4214 86522
rect 4266 86470 4278 86522
rect 4330 86470 4342 86522
rect 4394 86470 4406 86522
rect 4458 86470 4470 86522
rect 4522 86470 34934 86522
rect 34986 86470 34998 86522
rect 35050 86470 35062 86522
rect 35114 86470 35126 86522
rect 35178 86470 35190 86522
rect 35242 86470 65654 86522
rect 65706 86470 65718 86522
rect 65770 86470 65782 86522
rect 65834 86470 65846 86522
rect 65898 86470 65910 86522
rect 65962 86470 78844 86522
rect 1104 86448 78844 86470
rect 1397 86207 1455 86213
rect 1397 86173 1409 86207
rect 1443 86204 1455 86207
rect 2038 86204 2044 86216
rect 1443 86176 2044 86204
rect 1443 86173 1455 86176
rect 1397 86167 1455 86173
rect 2038 86164 2044 86176
rect 2096 86164 2102 86216
rect 1578 86068 1584 86080
rect 1539 86040 1584 86068
rect 1578 86028 1584 86040
rect 1636 86028 1642 86080
rect 1104 85978 78844 86000
rect 1104 85926 19574 85978
rect 19626 85926 19638 85978
rect 19690 85926 19702 85978
rect 19754 85926 19766 85978
rect 19818 85926 19830 85978
rect 19882 85926 50294 85978
rect 50346 85926 50358 85978
rect 50410 85926 50422 85978
rect 50474 85926 50486 85978
rect 50538 85926 50550 85978
rect 50602 85926 78844 85978
rect 1104 85904 78844 85926
rect 1104 85434 78844 85456
rect 1104 85382 4214 85434
rect 4266 85382 4278 85434
rect 4330 85382 4342 85434
rect 4394 85382 4406 85434
rect 4458 85382 4470 85434
rect 4522 85382 34934 85434
rect 34986 85382 34998 85434
rect 35050 85382 35062 85434
rect 35114 85382 35126 85434
rect 35178 85382 35190 85434
rect 35242 85382 65654 85434
rect 65706 85382 65718 85434
rect 65770 85382 65782 85434
rect 65834 85382 65846 85434
rect 65898 85382 65910 85434
rect 65962 85382 78844 85434
rect 1104 85360 78844 85382
rect 1104 84890 78844 84912
rect 1104 84838 19574 84890
rect 19626 84838 19638 84890
rect 19690 84838 19702 84890
rect 19754 84838 19766 84890
rect 19818 84838 19830 84890
rect 19882 84838 50294 84890
rect 50346 84838 50358 84890
rect 50410 84838 50422 84890
rect 50474 84838 50486 84890
rect 50538 84838 50550 84890
rect 50602 84838 78844 84890
rect 1104 84816 78844 84838
rect 1104 84346 78844 84368
rect 1104 84294 4214 84346
rect 4266 84294 4278 84346
rect 4330 84294 4342 84346
rect 4394 84294 4406 84346
rect 4458 84294 4470 84346
rect 4522 84294 34934 84346
rect 34986 84294 34998 84346
rect 35050 84294 35062 84346
rect 35114 84294 35126 84346
rect 35178 84294 35190 84346
rect 35242 84294 65654 84346
rect 65706 84294 65718 84346
rect 65770 84294 65782 84346
rect 65834 84294 65846 84346
rect 65898 84294 65910 84346
rect 65962 84294 78844 84346
rect 1104 84272 78844 84294
rect 1104 83802 78844 83824
rect 1104 83750 19574 83802
rect 19626 83750 19638 83802
rect 19690 83750 19702 83802
rect 19754 83750 19766 83802
rect 19818 83750 19830 83802
rect 19882 83750 50294 83802
rect 50346 83750 50358 83802
rect 50410 83750 50422 83802
rect 50474 83750 50486 83802
rect 50538 83750 50550 83802
rect 50602 83750 78844 83802
rect 1104 83728 78844 83750
rect 77662 83552 77668 83564
rect 77623 83524 77668 83552
rect 77662 83512 77668 83524
rect 77720 83512 77726 83564
rect 77846 83348 77852 83360
rect 77807 83320 77852 83348
rect 77846 83308 77852 83320
rect 77904 83308 77910 83360
rect 1104 83258 78844 83280
rect 1104 83206 4214 83258
rect 4266 83206 4278 83258
rect 4330 83206 4342 83258
rect 4394 83206 4406 83258
rect 4458 83206 4470 83258
rect 4522 83206 34934 83258
rect 34986 83206 34998 83258
rect 35050 83206 35062 83258
rect 35114 83206 35126 83258
rect 35178 83206 35190 83258
rect 35242 83206 65654 83258
rect 65706 83206 65718 83258
rect 65770 83206 65782 83258
rect 65834 83206 65846 83258
rect 65898 83206 65910 83258
rect 65962 83206 78844 83258
rect 1104 83184 78844 83206
rect 1104 82714 78844 82736
rect 1104 82662 19574 82714
rect 19626 82662 19638 82714
rect 19690 82662 19702 82714
rect 19754 82662 19766 82714
rect 19818 82662 19830 82714
rect 19882 82662 50294 82714
rect 50346 82662 50358 82714
rect 50410 82662 50422 82714
rect 50474 82662 50486 82714
rect 50538 82662 50550 82714
rect 50602 82662 78844 82714
rect 1104 82640 78844 82662
rect 1104 82170 78844 82192
rect 1104 82118 4214 82170
rect 4266 82118 4278 82170
rect 4330 82118 4342 82170
rect 4394 82118 4406 82170
rect 4458 82118 4470 82170
rect 4522 82118 34934 82170
rect 34986 82118 34998 82170
rect 35050 82118 35062 82170
rect 35114 82118 35126 82170
rect 35178 82118 35190 82170
rect 35242 82118 65654 82170
rect 65706 82118 65718 82170
rect 65770 82118 65782 82170
rect 65834 82118 65846 82170
rect 65898 82118 65910 82170
rect 65962 82118 78844 82170
rect 1104 82096 78844 82118
rect 1394 81852 1400 81864
rect 1355 81824 1400 81852
rect 1394 81812 1400 81824
rect 1452 81812 1458 81864
rect 1673 81787 1731 81793
rect 1673 81753 1685 81787
rect 1719 81784 1731 81787
rect 2130 81784 2136 81796
rect 1719 81756 2136 81784
rect 1719 81753 1731 81756
rect 1673 81747 1731 81753
rect 2130 81744 2136 81756
rect 2188 81744 2194 81796
rect 1104 81626 78844 81648
rect 1104 81574 19574 81626
rect 19626 81574 19638 81626
rect 19690 81574 19702 81626
rect 19754 81574 19766 81626
rect 19818 81574 19830 81626
rect 19882 81574 50294 81626
rect 50346 81574 50358 81626
rect 50410 81574 50422 81626
rect 50474 81574 50486 81626
rect 50538 81574 50550 81626
rect 50602 81574 78844 81626
rect 1104 81552 78844 81574
rect 1104 81082 78844 81104
rect 1104 81030 4214 81082
rect 4266 81030 4278 81082
rect 4330 81030 4342 81082
rect 4394 81030 4406 81082
rect 4458 81030 4470 81082
rect 4522 81030 34934 81082
rect 34986 81030 34998 81082
rect 35050 81030 35062 81082
rect 35114 81030 35126 81082
rect 35178 81030 35190 81082
rect 35242 81030 65654 81082
rect 65706 81030 65718 81082
rect 65770 81030 65782 81082
rect 65834 81030 65846 81082
rect 65898 81030 65910 81082
rect 65962 81030 78844 81082
rect 1104 81008 78844 81030
rect 1104 80538 78844 80560
rect 1104 80486 19574 80538
rect 19626 80486 19638 80538
rect 19690 80486 19702 80538
rect 19754 80486 19766 80538
rect 19818 80486 19830 80538
rect 19882 80486 50294 80538
rect 50346 80486 50358 80538
rect 50410 80486 50422 80538
rect 50474 80486 50486 80538
rect 50538 80486 50550 80538
rect 50602 80486 78844 80538
rect 1104 80464 78844 80486
rect 1104 79994 78844 80016
rect 1104 79942 4214 79994
rect 4266 79942 4278 79994
rect 4330 79942 4342 79994
rect 4394 79942 4406 79994
rect 4458 79942 4470 79994
rect 4522 79942 34934 79994
rect 34986 79942 34998 79994
rect 35050 79942 35062 79994
rect 35114 79942 35126 79994
rect 35178 79942 35190 79994
rect 35242 79942 65654 79994
rect 65706 79942 65718 79994
rect 65770 79942 65782 79994
rect 65834 79942 65846 79994
rect 65898 79942 65910 79994
rect 65962 79942 78844 79994
rect 1104 79920 78844 79942
rect 1104 79450 78844 79472
rect 1104 79398 19574 79450
rect 19626 79398 19638 79450
rect 19690 79398 19702 79450
rect 19754 79398 19766 79450
rect 19818 79398 19830 79450
rect 19882 79398 50294 79450
rect 50346 79398 50358 79450
rect 50410 79398 50422 79450
rect 50474 79398 50486 79450
rect 50538 79398 50550 79450
rect 50602 79398 78844 79450
rect 1104 79376 78844 79398
rect 10686 79336 10692 79348
rect 10647 79308 10692 79336
rect 10686 79296 10692 79308
rect 10744 79296 10750 79348
rect 2774 79160 2780 79212
rect 2832 79200 2838 79212
rect 10597 79203 10655 79209
rect 10597 79200 10609 79203
rect 2832 79172 10609 79200
rect 2832 79160 2838 79172
rect 10597 79169 10609 79172
rect 10643 79169 10655 79203
rect 77570 79200 77576 79212
rect 77531 79172 77576 79200
rect 10597 79163 10655 79169
rect 77570 79160 77576 79172
rect 77628 79160 77634 79212
rect 39942 78956 39948 79008
rect 40000 78996 40006 79008
rect 77665 78999 77723 79005
rect 77665 78996 77677 78999
rect 40000 78968 77677 78996
rect 40000 78956 40006 78968
rect 77665 78965 77677 78968
rect 77711 78965 77723 78999
rect 77665 78959 77723 78965
rect 1104 78906 78844 78928
rect 1104 78854 4214 78906
rect 4266 78854 4278 78906
rect 4330 78854 4342 78906
rect 4394 78854 4406 78906
rect 4458 78854 4470 78906
rect 4522 78854 34934 78906
rect 34986 78854 34998 78906
rect 35050 78854 35062 78906
rect 35114 78854 35126 78906
rect 35178 78854 35190 78906
rect 35242 78854 65654 78906
rect 65706 78854 65718 78906
rect 65770 78854 65782 78906
rect 65834 78854 65846 78906
rect 65898 78854 65910 78906
rect 65962 78854 78844 78906
rect 1104 78832 78844 78854
rect 1397 78591 1455 78597
rect 1397 78557 1409 78591
rect 1443 78588 1455 78591
rect 2590 78588 2596 78600
rect 1443 78560 2596 78588
rect 1443 78557 1455 78560
rect 1397 78551 1455 78557
rect 2590 78548 2596 78560
rect 2648 78548 2654 78600
rect 1578 78452 1584 78464
rect 1539 78424 1584 78452
rect 1578 78412 1584 78424
rect 1636 78412 1642 78464
rect 1104 78362 78844 78384
rect 1104 78310 19574 78362
rect 19626 78310 19638 78362
rect 19690 78310 19702 78362
rect 19754 78310 19766 78362
rect 19818 78310 19830 78362
rect 19882 78310 50294 78362
rect 50346 78310 50358 78362
rect 50410 78310 50422 78362
rect 50474 78310 50486 78362
rect 50538 78310 50550 78362
rect 50602 78310 78844 78362
rect 1104 78288 78844 78310
rect 2590 78248 2596 78260
rect 2551 78220 2596 78248
rect 2590 78208 2596 78220
rect 2648 78208 2654 78260
rect 2774 78112 2780 78124
rect 2735 78084 2780 78112
rect 2774 78072 2780 78084
rect 2832 78112 2838 78124
rect 3050 78112 3056 78124
rect 2832 78084 3056 78112
rect 2832 78072 2838 78084
rect 3050 78072 3056 78084
rect 3108 78072 3114 78124
rect 1104 77818 78844 77840
rect 1104 77766 4214 77818
rect 4266 77766 4278 77818
rect 4330 77766 4342 77818
rect 4394 77766 4406 77818
rect 4458 77766 4470 77818
rect 4522 77766 34934 77818
rect 34986 77766 34998 77818
rect 35050 77766 35062 77818
rect 35114 77766 35126 77818
rect 35178 77766 35190 77818
rect 35242 77766 65654 77818
rect 65706 77766 65718 77818
rect 65770 77766 65782 77818
rect 65834 77766 65846 77818
rect 65898 77766 65910 77818
rect 65962 77766 78844 77818
rect 1104 77744 78844 77766
rect 1104 77274 78844 77296
rect 1104 77222 19574 77274
rect 19626 77222 19638 77274
rect 19690 77222 19702 77274
rect 19754 77222 19766 77274
rect 19818 77222 19830 77274
rect 19882 77222 50294 77274
rect 50346 77222 50358 77274
rect 50410 77222 50422 77274
rect 50474 77222 50486 77274
rect 50538 77222 50550 77274
rect 50602 77222 78844 77274
rect 1104 77200 78844 77222
rect 1104 76730 78844 76752
rect 1104 76678 4214 76730
rect 4266 76678 4278 76730
rect 4330 76678 4342 76730
rect 4394 76678 4406 76730
rect 4458 76678 4470 76730
rect 4522 76678 34934 76730
rect 34986 76678 34998 76730
rect 35050 76678 35062 76730
rect 35114 76678 35126 76730
rect 35178 76678 35190 76730
rect 35242 76678 65654 76730
rect 65706 76678 65718 76730
rect 65770 76678 65782 76730
rect 65834 76678 65846 76730
rect 65898 76678 65910 76730
rect 65962 76678 78844 76730
rect 1104 76656 78844 76678
rect 1104 76186 78844 76208
rect 1104 76134 19574 76186
rect 19626 76134 19638 76186
rect 19690 76134 19702 76186
rect 19754 76134 19766 76186
rect 19818 76134 19830 76186
rect 19882 76134 50294 76186
rect 50346 76134 50358 76186
rect 50410 76134 50422 76186
rect 50474 76134 50486 76186
rect 50538 76134 50550 76186
rect 50602 76134 78844 76186
rect 1104 76112 78844 76134
rect 1104 75642 78844 75664
rect 1104 75590 4214 75642
rect 4266 75590 4278 75642
rect 4330 75590 4342 75642
rect 4394 75590 4406 75642
rect 4458 75590 4470 75642
rect 4522 75590 34934 75642
rect 34986 75590 34998 75642
rect 35050 75590 35062 75642
rect 35114 75590 35126 75642
rect 35178 75590 35190 75642
rect 35242 75590 65654 75642
rect 65706 75590 65718 75642
rect 65770 75590 65782 75642
rect 65834 75590 65846 75642
rect 65898 75590 65910 75642
rect 65962 75590 78844 75642
rect 1104 75568 78844 75590
rect 77849 75327 77907 75333
rect 77849 75293 77861 75327
rect 77895 75324 77907 75327
rect 77938 75324 77944 75336
rect 77895 75296 77944 75324
rect 77895 75293 77907 75296
rect 77849 75287 77907 75293
rect 77938 75284 77944 75296
rect 77996 75284 78002 75336
rect 78030 75188 78036 75200
rect 77991 75160 78036 75188
rect 78030 75148 78036 75160
rect 78088 75148 78094 75200
rect 1104 75098 78844 75120
rect 1104 75046 19574 75098
rect 19626 75046 19638 75098
rect 19690 75046 19702 75098
rect 19754 75046 19766 75098
rect 19818 75046 19830 75098
rect 19882 75046 50294 75098
rect 50346 75046 50358 75098
rect 50410 75046 50422 75098
rect 50474 75046 50486 75098
rect 50538 75046 50550 75098
rect 50602 75046 78844 75098
rect 1104 75024 78844 75046
rect 1104 74554 78844 74576
rect 1104 74502 4214 74554
rect 4266 74502 4278 74554
rect 4330 74502 4342 74554
rect 4394 74502 4406 74554
rect 4458 74502 4470 74554
rect 4522 74502 34934 74554
rect 34986 74502 34998 74554
rect 35050 74502 35062 74554
rect 35114 74502 35126 74554
rect 35178 74502 35190 74554
rect 35242 74502 65654 74554
rect 65706 74502 65718 74554
rect 65770 74502 65782 74554
rect 65834 74502 65846 74554
rect 65898 74502 65910 74554
rect 65962 74502 78844 74554
rect 1104 74480 78844 74502
rect 1670 74264 1676 74316
rect 1728 74304 1734 74316
rect 1946 74304 1952 74316
rect 1728 74276 1952 74304
rect 1728 74264 1734 74276
rect 1946 74264 1952 74276
rect 2004 74264 2010 74316
rect 1397 74239 1455 74245
rect 1397 74205 1409 74239
rect 1443 74236 1455 74239
rect 1486 74236 1492 74248
rect 1443 74208 1492 74236
rect 1443 74205 1455 74208
rect 1397 74199 1455 74205
rect 1486 74196 1492 74208
rect 1544 74196 1550 74248
rect 1578 74100 1584 74112
rect 1539 74072 1584 74100
rect 1578 74060 1584 74072
rect 1636 74060 1642 74112
rect 1104 74010 78844 74032
rect 1104 73958 19574 74010
rect 19626 73958 19638 74010
rect 19690 73958 19702 74010
rect 19754 73958 19766 74010
rect 19818 73958 19830 74010
rect 19882 73958 50294 74010
rect 50346 73958 50358 74010
rect 50410 73958 50422 74010
rect 50474 73958 50486 74010
rect 50538 73958 50550 74010
rect 50602 73958 78844 74010
rect 1104 73936 78844 73958
rect 1104 73466 78844 73488
rect 1104 73414 4214 73466
rect 4266 73414 4278 73466
rect 4330 73414 4342 73466
rect 4394 73414 4406 73466
rect 4458 73414 4470 73466
rect 4522 73414 34934 73466
rect 34986 73414 34998 73466
rect 35050 73414 35062 73466
rect 35114 73414 35126 73466
rect 35178 73414 35190 73466
rect 35242 73414 65654 73466
rect 65706 73414 65718 73466
rect 65770 73414 65782 73466
rect 65834 73414 65846 73466
rect 65898 73414 65910 73466
rect 65962 73414 78844 73466
rect 1104 73392 78844 73414
rect 1104 72922 78844 72944
rect 1104 72870 19574 72922
rect 19626 72870 19638 72922
rect 19690 72870 19702 72922
rect 19754 72870 19766 72922
rect 19818 72870 19830 72922
rect 19882 72870 50294 72922
rect 50346 72870 50358 72922
rect 50410 72870 50422 72922
rect 50474 72870 50486 72922
rect 50538 72870 50550 72922
rect 50602 72870 78844 72922
rect 1104 72848 78844 72870
rect 1104 72378 78844 72400
rect 1104 72326 4214 72378
rect 4266 72326 4278 72378
rect 4330 72326 4342 72378
rect 4394 72326 4406 72378
rect 4458 72326 4470 72378
rect 4522 72326 34934 72378
rect 34986 72326 34998 72378
rect 35050 72326 35062 72378
rect 35114 72326 35126 72378
rect 35178 72326 35190 72378
rect 35242 72326 65654 72378
rect 65706 72326 65718 72378
rect 65770 72326 65782 72378
rect 65834 72326 65846 72378
rect 65898 72326 65910 72378
rect 65962 72326 78844 72378
rect 1104 72304 78844 72326
rect 67821 72063 67879 72069
rect 67821 72029 67833 72063
rect 67867 72060 67879 72063
rect 76742 72060 76748 72072
rect 67867 72032 76748 72060
rect 67867 72029 67879 72032
rect 67821 72023 67879 72029
rect 76742 72020 76748 72032
rect 76800 72020 76806 72072
rect 45186 71952 45192 72004
rect 45244 71992 45250 72004
rect 68097 71995 68155 72001
rect 68097 71992 68109 71995
rect 45244 71964 68109 71992
rect 45244 71952 45250 71964
rect 68097 71961 68109 71964
rect 68143 71961 68155 71995
rect 68097 71955 68155 71961
rect 1104 71834 78844 71856
rect 1104 71782 19574 71834
rect 19626 71782 19638 71834
rect 19690 71782 19702 71834
rect 19754 71782 19766 71834
rect 19818 71782 19830 71834
rect 19882 71782 50294 71834
rect 50346 71782 50358 71834
rect 50410 71782 50422 71834
rect 50474 71782 50486 71834
rect 50538 71782 50550 71834
rect 50602 71782 78844 71834
rect 1104 71760 78844 71782
rect 76558 71544 76564 71596
rect 76616 71584 76622 71596
rect 77665 71587 77723 71593
rect 77665 71584 77677 71587
rect 76616 71556 77677 71584
rect 76616 71544 76622 71556
rect 77665 71553 77677 71556
rect 77711 71553 77723 71587
rect 77665 71547 77723 71553
rect 77846 71448 77852 71460
rect 77807 71420 77852 71448
rect 77846 71408 77852 71420
rect 77904 71408 77910 71460
rect 1104 71290 78844 71312
rect 1104 71238 4214 71290
rect 4266 71238 4278 71290
rect 4330 71238 4342 71290
rect 4394 71238 4406 71290
rect 4458 71238 4470 71290
rect 4522 71238 34934 71290
rect 34986 71238 34998 71290
rect 35050 71238 35062 71290
rect 35114 71238 35126 71290
rect 35178 71238 35190 71290
rect 35242 71238 65654 71290
rect 65706 71238 65718 71290
rect 65770 71238 65782 71290
rect 65834 71238 65846 71290
rect 65898 71238 65910 71290
rect 65962 71238 78844 71290
rect 1104 71216 78844 71238
rect 76558 71176 76564 71188
rect 76519 71148 76564 71176
rect 76558 71136 76564 71148
rect 76616 71136 76622 71188
rect 2038 71108 2044 71120
rect 1999 71080 2044 71108
rect 2038 71068 2044 71080
rect 2096 71068 2102 71120
rect 76742 70972 76748 70984
rect 76655 70944 76748 70972
rect 76742 70932 76748 70944
rect 76800 70972 76806 70984
rect 77662 70972 77668 70984
rect 76800 70944 77668 70972
rect 76800 70932 76806 70944
rect 77662 70932 77668 70944
rect 77720 70932 77726 70984
rect 1670 70864 1676 70916
rect 1728 70904 1734 70916
rect 1857 70907 1915 70913
rect 1857 70904 1869 70907
rect 1728 70876 1869 70904
rect 1728 70864 1734 70876
rect 1857 70873 1869 70876
rect 1903 70873 1915 70907
rect 1857 70867 1915 70873
rect 1104 70746 78844 70768
rect 1104 70694 19574 70746
rect 19626 70694 19638 70746
rect 19690 70694 19702 70746
rect 19754 70694 19766 70746
rect 19818 70694 19830 70746
rect 19882 70694 50294 70746
rect 50346 70694 50358 70746
rect 50410 70694 50422 70746
rect 50474 70694 50486 70746
rect 50538 70694 50550 70746
rect 50602 70694 78844 70746
rect 1104 70672 78844 70694
rect 1394 70496 1400 70508
rect 1355 70468 1400 70496
rect 1394 70456 1400 70468
rect 1452 70456 1458 70508
rect 1578 70292 1584 70304
rect 1539 70264 1584 70292
rect 1578 70252 1584 70264
rect 1636 70252 1642 70304
rect 1104 70202 78844 70224
rect 1104 70150 4214 70202
rect 4266 70150 4278 70202
rect 4330 70150 4342 70202
rect 4394 70150 4406 70202
rect 4458 70150 4470 70202
rect 4522 70150 34934 70202
rect 34986 70150 34998 70202
rect 35050 70150 35062 70202
rect 35114 70150 35126 70202
rect 35178 70150 35190 70202
rect 35242 70150 65654 70202
rect 65706 70150 65718 70202
rect 65770 70150 65782 70202
rect 65834 70150 65846 70202
rect 65898 70150 65910 70202
rect 65962 70150 78844 70202
rect 1104 70128 78844 70150
rect 1394 70048 1400 70100
rect 1452 70088 1458 70100
rect 1765 70091 1823 70097
rect 1765 70088 1777 70091
rect 1452 70060 1777 70088
rect 1452 70048 1458 70060
rect 1765 70057 1777 70060
rect 1811 70057 1823 70091
rect 1765 70051 1823 70057
rect 1670 69844 1676 69896
rect 1728 69884 1734 69896
rect 1949 69887 2007 69893
rect 1949 69884 1961 69887
rect 1728 69856 1961 69884
rect 1728 69844 1734 69856
rect 1949 69853 1961 69856
rect 1995 69853 2007 69887
rect 1949 69847 2007 69853
rect 77478 69708 77484 69760
rect 77536 69748 77542 69760
rect 77938 69748 77944 69760
rect 77536 69720 77944 69748
rect 77536 69708 77542 69720
rect 77938 69708 77944 69720
rect 77996 69708 78002 69760
rect 1104 69658 78844 69680
rect 1104 69606 19574 69658
rect 19626 69606 19638 69658
rect 19690 69606 19702 69658
rect 19754 69606 19766 69658
rect 19818 69606 19830 69658
rect 19882 69606 50294 69658
rect 50346 69606 50358 69658
rect 50410 69606 50422 69658
rect 50474 69606 50486 69658
rect 50538 69606 50550 69658
rect 50602 69606 78844 69658
rect 1104 69584 78844 69606
rect 1104 69114 78844 69136
rect 1104 69062 4214 69114
rect 4266 69062 4278 69114
rect 4330 69062 4342 69114
rect 4394 69062 4406 69114
rect 4458 69062 4470 69114
rect 4522 69062 34934 69114
rect 34986 69062 34998 69114
rect 35050 69062 35062 69114
rect 35114 69062 35126 69114
rect 35178 69062 35190 69114
rect 35242 69062 65654 69114
rect 65706 69062 65718 69114
rect 65770 69062 65782 69114
rect 65834 69062 65846 69114
rect 65898 69062 65910 69114
rect 65962 69062 78844 69114
rect 1104 69040 78844 69062
rect 1104 68570 78844 68592
rect 1104 68518 19574 68570
rect 19626 68518 19638 68570
rect 19690 68518 19702 68570
rect 19754 68518 19766 68570
rect 19818 68518 19830 68570
rect 19882 68518 50294 68570
rect 50346 68518 50358 68570
rect 50410 68518 50422 68570
rect 50474 68518 50486 68570
rect 50538 68518 50550 68570
rect 50602 68518 78844 68570
rect 1104 68496 78844 68518
rect 1104 68026 78844 68048
rect 1104 67974 4214 68026
rect 4266 67974 4278 68026
rect 4330 67974 4342 68026
rect 4394 67974 4406 68026
rect 4458 67974 4470 68026
rect 4522 67974 34934 68026
rect 34986 67974 34998 68026
rect 35050 67974 35062 68026
rect 35114 67974 35126 68026
rect 35178 67974 35190 68026
rect 35242 67974 65654 68026
rect 65706 67974 65718 68026
rect 65770 67974 65782 68026
rect 65834 67974 65846 68026
rect 65898 67974 65910 68026
rect 65962 67974 78844 68026
rect 1104 67952 78844 67974
rect 77757 67643 77815 67649
rect 77757 67609 77769 67643
rect 77803 67640 77815 67643
rect 77938 67640 77944 67652
rect 77803 67612 77944 67640
rect 77803 67609 77815 67612
rect 77757 67603 77815 67609
rect 77938 67600 77944 67612
rect 77996 67600 78002 67652
rect 77846 67572 77852 67584
rect 77807 67544 77852 67572
rect 77846 67532 77852 67544
rect 77904 67532 77910 67584
rect 1104 67482 78844 67504
rect 1104 67430 19574 67482
rect 19626 67430 19638 67482
rect 19690 67430 19702 67482
rect 19754 67430 19766 67482
rect 19818 67430 19830 67482
rect 19882 67430 50294 67482
rect 50346 67430 50358 67482
rect 50410 67430 50422 67482
rect 50474 67430 50486 67482
rect 50538 67430 50550 67482
rect 50602 67430 78844 67482
rect 1104 67408 78844 67430
rect 1104 66938 78844 66960
rect 1104 66886 4214 66938
rect 4266 66886 4278 66938
rect 4330 66886 4342 66938
rect 4394 66886 4406 66938
rect 4458 66886 4470 66938
rect 4522 66886 34934 66938
rect 34986 66886 34998 66938
rect 35050 66886 35062 66938
rect 35114 66886 35126 66938
rect 35178 66886 35190 66938
rect 35242 66886 65654 66938
rect 65706 66886 65718 66938
rect 65770 66886 65782 66938
rect 65834 66886 65846 66938
rect 65898 66886 65910 66938
rect 65962 66886 78844 66938
rect 1104 66864 78844 66886
rect 1104 66394 78844 66416
rect 1104 66342 19574 66394
rect 19626 66342 19638 66394
rect 19690 66342 19702 66394
rect 19754 66342 19766 66394
rect 19818 66342 19830 66394
rect 19882 66342 50294 66394
rect 50346 66342 50358 66394
rect 50410 66342 50422 66394
rect 50474 66342 50486 66394
rect 50538 66342 50550 66394
rect 50602 66342 78844 66394
rect 1104 66320 78844 66342
rect 1397 66147 1455 66153
rect 1397 66113 1409 66147
rect 1443 66144 1455 66147
rect 2314 66144 2320 66156
rect 1443 66116 2176 66144
rect 2275 66116 2320 66144
rect 1443 66113 1455 66116
rect 1397 66107 1455 66113
rect 1578 66008 1584 66020
rect 1539 65980 1584 66008
rect 1578 65968 1584 65980
rect 1636 65968 1642 66020
rect 2148 66017 2176 66116
rect 2314 66104 2320 66116
rect 2372 66104 2378 66156
rect 2133 66011 2191 66017
rect 2133 65977 2145 66011
rect 2179 65977 2191 66011
rect 2133 65971 2191 65977
rect 1104 65850 78844 65872
rect 1104 65798 4214 65850
rect 4266 65798 4278 65850
rect 4330 65798 4342 65850
rect 4394 65798 4406 65850
rect 4458 65798 4470 65850
rect 4522 65798 34934 65850
rect 34986 65798 34998 65850
rect 35050 65798 35062 65850
rect 35114 65798 35126 65850
rect 35178 65798 35190 65850
rect 35242 65798 65654 65850
rect 65706 65798 65718 65850
rect 65770 65798 65782 65850
rect 65834 65798 65846 65850
rect 65898 65798 65910 65850
rect 65962 65798 78844 65850
rect 1104 65776 78844 65798
rect 40678 65560 40684 65612
rect 40736 65600 40742 65612
rect 41877 65603 41935 65609
rect 41877 65600 41889 65603
rect 40736 65572 41889 65600
rect 40736 65560 40742 65572
rect 41877 65569 41889 65572
rect 41923 65569 41935 65603
rect 41877 65563 41935 65569
rect 1857 65535 1915 65541
rect 1857 65501 1869 65535
rect 1903 65532 1915 65535
rect 2314 65532 2320 65544
rect 1903 65504 2320 65532
rect 1903 65501 1915 65504
rect 1857 65495 1915 65501
rect 2314 65492 2320 65504
rect 2372 65492 2378 65544
rect 39850 65532 39856 65544
rect 39811 65504 39856 65532
rect 39850 65492 39856 65504
rect 39908 65492 39914 65544
rect 11882 65424 11888 65476
rect 11940 65464 11946 65476
rect 11940 65436 26234 65464
rect 11940 65424 11946 65436
rect 1762 65356 1768 65408
rect 1820 65396 1826 65408
rect 1949 65399 2007 65405
rect 1949 65396 1961 65399
rect 1820 65368 1961 65396
rect 1820 65356 1826 65368
rect 1949 65365 1961 65368
rect 1995 65365 2007 65399
rect 26206 65396 26234 65436
rect 40034 65424 40040 65476
rect 40092 65464 40098 65476
rect 40129 65467 40187 65473
rect 40129 65464 40141 65467
rect 40092 65436 40141 65464
rect 40092 65424 40098 65436
rect 40129 65433 40141 65436
rect 40175 65433 40187 65467
rect 40129 65427 40187 65433
rect 40236 65436 40618 65464
rect 40236 65396 40264 65436
rect 26206 65368 40264 65396
rect 1949 65359 2007 65365
rect 1104 65306 78844 65328
rect 1104 65254 19574 65306
rect 19626 65254 19638 65306
rect 19690 65254 19702 65306
rect 19754 65254 19766 65306
rect 19818 65254 19830 65306
rect 19882 65254 50294 65306
rect 50346 65254 50358 65306
rect 50410 65254 50422 65306
rect 50474 65254 50486 65306
rect 50538 65254 50550 65306
rect 50602 65254 78844 65306
rect 1104 65232 78844 65254
rect 40034 65192 40040 65204
rect 39995 65164 40040 65192
rect 40034 65152 40040 65164
rect 40092 65152 40098 65204
rect 41046 65192 41052 65204
rect 41007 65164 41052 65192
rect 41046 65152 41052 65164
rect 41104 65152 41110 65204
rect 40221 65059 40279 65065
rect 40221 65025 40233 65059
rect 40267 65056 40279 65059
rect 40267 65028 41276 65056
rect 40267 65025 40279 65028
rect 40221 65019 40279 65025
rect 40678 64988 40684 65000
rect 40639 64960 40684 64988
rect 40678 64948 40684 64960
rect 40736 64948 40742 65000
rect 41248 64929 41276 65028
rect 41233 64923 41291 64929
rect 41233 64889 41245 64923
rect 41279 64889 41291 64923
rect 41233 64883 41291 64889
rect 40862 64812 40868 64864
rect 40920 64852 40926 64864
rect 41049 64855 41107 64861
rect 41049 64852 41061 64855
rect 40920 64824 41061 64852
rect 40920 64812 40926 64824
rect 41049 64821 41061 64824
rect 41095 64821 41107 64855
rect 41049 64815 41107 64821
rect 41690 64812 41696 64864
rect 41748 64852 41754 64864
rect 77846 64852 77852 64864
rect 41748 64824 77852 64852
rect 41748 64812 41754 64824
rect 77846 64812 77852 64824
rect 77904 64812 77910 64864
rect 1104 64762 78844 64784
rect 1104 64710 4214 64762
rect 4266 64710 4278 64762
rect 4330 64710 4342 64762
rect 4394 64710 4406 64762
rect 4458 64710 4470 64762
rect 4522 64710 34934 64762
rect 34986 64710 34998 64762
rect 35050 64710 35062 64762
rect 35114 64710 35126 64762
rect 35178 64710 35190 64762
rect 35242 64710 65654 64762
rect 65706 64710 65718 64762
rect 65770 64710 65782 64762
rect 65834 64710 65846 64762
rect 65898 64710 65910 64762
rect 65962 64710 78844 64762
rect 1104 64688 78844 64710
rect 41690 64580 41696 64592
rect 40052 64552 41696 64580
rect 39482 64404 39488 64456
rect 39540 64444 39546 64456
rect 40052 64453 40080 64552
rect 41690 64540 41696 64552
rect 41748 64540 41754 64592
rect 41046 64512 41052 64524
rect 40788 64484 41052 64512
rect 40037 64447 40095 64453
rect 40037 64444 40049 64447
rect 39540 64416 40049 64444
rect 39540 64404 39546 64416
rect 40037 64413 40049 64416
rect 40083 64413 40095 64447
rect 40494 64444 40500 64456
rect 40455 64416 40500 64444
rect 40037 64407 40095 64413
rect 40494 64404 40500 64416
rect 40552 64404 40558 64456
rect 40788 64453 40816 64484
rect 41046 64472 41052 64484
rect 41104 64472 41110 64524
rect 40773 64447 40831 64453
rect 40773 64413 40785 64447
rect 40819 64413 40831 64447
rect 40773 64407 40831 64413
rect 40862 64404 40868 64456
rect 40920 64444 40926 64456
rect 40920 64416 40965 64444
rect 40920 64404 40926 64416
rect 1104 64218 78844 64240
rect 1104 64166 19574 64218
rect 19626 64166 19638 64218
rect 19690 64166 19702 64218
rect 19754 64166 19766 64218
rect 19818 64166 19830 64218
rect 19882 64166 50294 64218
rect 50346 64166 50358 64218
rect 50410 64166 50422 64218
rect 50474 64166 50486 64218
rect 50538 64166 50550 64218
rect 50602 64166 78844 64218
rect 1104 64144 78844 64166
rect 39482 63968 39488 63980
rect 39443 63940 39488 63968
rect 39482 63928 39488 63940
rect 39540 63928 39546 63980
rect 39482 63724 39488 63776
rect 39540 63764 39546 63776
rect 39577 63767 39635 63773
rect 39577 63764 39589 63767
rect 39540 63736 39589 63764
rect 39540 63724 39546 63736
rect 39577 63733 39589 63736
rect 39623 63733 39635 63767
rect 39577 63727 39635 63733
rect 1104 63674 78844 63696
rect 1104 63622 4214 63674
rect 4266 63622 4278 63674
rect 4330 63622 4342 63674
rect 4394 63622 4406 63674
rect 4458 63622 4470 63674
rect 4522 63622 34934 63674
rect 34986 63622 34998 63674
rect 35050 63622 35062 63674
rect 35114 63622 35126 63674
rect 35178 63622 35190 63674
rect 35242 63622 65654 63674
rect 65706 63622 65718 63674
rect 65770 63622 65782 63674
rect 65834 63622 65846 63674
rect 65898 63622 65910 63674
rect 65962 63622 78844 63674
rect 1104 63600 78844 63622
rect 38286 63316 38292 63368
rect 38344 63356 38350 63368
rect 77481 63359 77539 63365
rect 77481 63356 77493 63359
rect 38344 63328 77493 63356
rect 38344 63316 38350 63328
rect 77481 63325 77493 63328
rect 77527 63356 77539 63359
rect 77849 63359 77907 63365
rect 77849 63356 77861 63359
rect 77527 63328 77861 63356
rect 77527 63325 77539 63328
rect 77481 63319 77539 63325
rect 77849 63325 77861 63328
rect 77895 63325 77907 63359
rect 77849 63319 77907 63325
rect 78030 63220 78036 63232
rect 77991 63192 78036 63220
rect 78030 63180 78036 63192
rect 78088 63180 78094 63232
rect 1104 63130 78844 63152
rect 1104 63078 19574 63130
rect 19626 63078 19638 63130
rect 19690 63078 19702 63130
rect 19754 63078 19766 63130
rect 19818 63078 19830 63130
rect 19882 63078 50294 63130
rect 50346 63078 50358 63130
rect 50410 63078 50422 63130
rect 50474 63078 50486 63130
rect 50538 63078 50550 63130
rect 50602 63078 78844 63130
rect 1104 63056 78844 63078
rect 1394 62880 1400 62892
rect 1355 62852 1400 62880
rect 1394 62840 1400 62852
rect 1452 62840 1458 62892
rect 1578 62676 1584 62688
rect 1539 62648 1584 62676
rect 1578 62636 1584 62648
rect 1636 62636 1642 62688
rect 1104 62586 78844 62608
rect 1104 62534 4214 62586
rect 4266 62534 4278 62586
rect 4330 62534 4342 62586
rect 4394 62534 4406 62586
rect 4458 62534 4470 62586
rect 4522 62534 34934 62586
rect 34986 62534 34998 62586
rect 35050 62534 35062 62586
rect 35114 62534 35126 62586
rect 35178 62534 35190 62586
rect 35242 62534 65654 62586
rect 65706 62534 65718 62586
rect 65770 62534 65782 62586
rect 65834 62534 65846 62586
rect 65898 62534 65910 62586
rect 65962 62534 78844 62586
rect 1104 62512 78844 62534
rect 1104 62042 78844 62064
rect 1104 61990 19574 62042
rect 19626 61990 19638 62042
rect 19690 61990 19702 62042
rect 19754 61990 19766 62042
rect 19818 61990 19830 62042
rect 19882 61990 50294 62042
rect 50346 61990 50358 62042
rect 50410 61990 50422 62042
rect 50474 61990 50486 62042
rect 50538 61990 50550 62042
rect 50602 61990 78844 62042
rect 1104 61968 78844 61990
rect 1104 61498 78844 61520
rect 1104 61446 4214 61498
rect 4266 61446 4278 61498
rect 4330 61446 4342 61498
rect 4394 61446 4406 61498
rect 4458 61446 4470 61498
rect 4522 61446 34934 61498
rect 34986 61446 34998 61498
rect 35050 61446 35062 61498
rect 35114 61446 35126 61498
rect 35178 61446 35190 61498
rect 35242 61446 65654 61498
rect 65706 61446 65718 61498
rect 65770 61446 65782 61498
rect 65834 61446 65846 61498
rect 65898 61446 65910 61498
rect 65962 61446 78844 61498
rect 1104 61424 78844 61446
rect 39758 61140 39764 61192
rect 39816 61180 39822 61192
rect 39853 61183 39911 61189
rect 39853 61180 39865 61183
rect 39816 61152 39865 61180
rect 39816 61140 39822 61152
rect 39853 61149 39865 61152
rect 39899 61149 39911 61183
rect 39853 61143 39911 61149
rect 19426 61072 19432 61124
rect 19484 61112 19490 61124
rect 40129 61115 40187 61121
rect 40129 61112 40141 61115
rect 19484 61084 40141 61112
rect 19484 61072 19490 61084
rect 40129 61081 40141 61084
rect 40175 61081 40187 61115
rect 40129 61075 40187 61081
rect 1104 60954 78844 60976
rect 1104 60902 19574 60954
rect 19626 60902 19638 60954
rect 19690 60902 19702 60954
rect 19754 60902 19766 60954
rect 19818 60902 19830 60954
rect 19882 60902 50294 60954
rect 50346 60902 50358 60954
rect 50410 60902 50422 60954
rect 50474 60902 50486 60954
rect 50538 60902 50550 60954
rect 50602 60902 78844 60954
rect 1104 60880 78844 60902
rect 39942 60772 39948 60784
rect 39903 60744 39948 60772
rect 39942 60732 39948 60744
rect 40000 60732 40006 60784
rect 40770 60732 40776 60784
rect 40828 60772 40834 60784
rect 40865 60775 40923 60781
rect 40865 60772 40877 60775
rect 40828 60744 40877 60772
rect 40828 60732 40834 60744
rect 40865 60741 40877 60744
rect 40911 60741 40923 60775
rect 40865 60735 40923 60741
rect 38838 60664 38844 60716
rect 38896 60704 38902 60716
rect 38933 60707 38991 60713
rect 38933 60704 38945 60707
rect 38896 60676 38945 60704
rect 38896 60664 38902 60676
rect 38933 60673 38945 60676
rect 38979 60673 38991 60707
rect 38933 60667 38991 60673
rect 39209 60639 39267 60645
rect 39209 60605 39221 60639
rect 39255 60636 39267 60639
rect 77294 60636 77300 60648
rect 39255 60608 77300 60636
rect 39255 60605 39267 60608
rect 39209 60599 39267 60605
rect 77294 60596 77300 60608
rect 77352 60596 77358 60648
rect 1486 60528 1492 60580
rect 1544 60568 1550 60580
rect 40129 60571 40187 60577
rect 40129 60568 40141 60571
rect 1544 60540 40141 60568
rect 1544 60528 1550 60540
rect 40129 60537 40141 60540
rect 40175 60537 40187 60571
rect 40129 60531 40187 60537
rect 41141 60503 41199 60509
rect 41141 60469 41153 60503
rect 41187 60500 41199 60503
rect 77570 60500 77576 60512
rect 41187 60472 77576 60500
rect 41187 60469 41199 60472
rect 41141 60463 41199 60469
rect 77570 60460 77576 60472
rect 77628 60460 77634 60512
rect 1104 60410 78844 60432
rect 1104 60358 4214 60410
rect 4266 60358 4278 60410
rect 4330 60358 4342 60410
rect 4394 60358 4406 60410
rect 4458 60358 4470 60410
rect 4522 60358 34934 60410
rect 34986 60358 34998 60410
rect 35050 60358 35062 60410
rect 35114 60358 35126 60410
rect 35178 60358 35190 60410
rect 35242 60358 65654 60410
rect 65706 60358 65718 60410
rect 65770 60358 65782 60410
rect 65834 60358 65846 60410
rect 65898 60358 65910 60410
rect 65962 60358 78844 60410
rect 1104 60336 78844 60358
rect 2130 60256 2136 60308
rect 2188 60296 2194 60308
rect 35802 60296 35808 60308
rect 2188 60268 9674 60296
rect 35763 60268 35808 60296
rect 2188 60256 2194 60268
rect 1854 60120 1860 60172
rect 1912 60160 1918 60172
rect 9646 60160 9674 60268
rect 35802 60256 35808 60268
rect 35860 60256 35866 60308
rect 36354 60296 36360 60308
rect 36315 60268 36360 60296
rect 36354 60256 36360 60268
rect 36412 60256 36418 60308
rect 38286 60296 38292 60308
rect 38247 60268 38292 60296
rect 38286 60256 38292 60268
rect 38344 60256 38350 60308
rect 77754 60256 77760 60308
rect 77812 60296 77818 60308
rect 77849 60299 77907 60305
rect 77849 60296 77861 60299
rect 77812 60268 77861 60296
rect 77812 60256 77818 60268
rect 77849 60265 77861 60268
rect 77895 60265 77907 60299
rect 77849 60259 77907 60265
rect 26206 60200 41276 60228
rect 1912 60132 2360 60160
rect 9646 60132 21404 60160
rect 1912 60120 1918 60132
rect 1765 60095 1823 60101
rect 1765 60061 1777 60095
rect 1811 60092 1823 60095
rect 2222 60092 2228 60104
rect 1811 60064 2228 60092
rect 1811 60061 1823 60064
rect 1765 60055 1823 60061
rect 2222 60052 2228 60064
rect 2280 60052 2286 60104
rect 2332 60092 2360 60132
rect 19245 60095 19303 60101
rect 19245 60092 19257 60095
rect 2332 60064 19257 60092
rect 19245 60061 19257 60064
rect 19291 60061 19303 60095
rect 21376 60092 21404 60132
rect 22646 60120 22652 60172
rect 22704 60160 22710 60172
rect 26206 60160 26234 60200
rect 41248 60169 41276 60200
rect 41233 60163 41291 60169
rect 22704 60132 26234 60160
rect 37936 60132 39988 60160
rect 22704 60120 22710 60132
rect 37936 60092 37964 60132
rect 39960 60101 39988 60132
rect 41233 60129 41245 60163
rect 41279 60129 41291 60163
rect 41233 60123 41291 60129
rect 21376 60064 37964 60092
rect 38105 60095 38163 60101
rect 19245 60055 19303 60061
rect 38105 60061 38117 60095
rect 38151 60061 38163 60095
rect 38105 60055 38163 60061
rect 39945 60095 40003 60101
rect 39945 60061 39957 60095
rect 39991 60061 40003 60095
rect 41046 60092 41052 60104
rect 41007 60064 41052 60092
rect 39945 60055 40003 60061
rect 19521 60027 19579 60033
rect 19521 59993 19533 60027
rect 19567 60024 19579 60027
rect 19978 60024 19984 60036
rect 19567 59996 19984 60024
rect 19567 59993 19579 59996
rect 19521 59987 19579 59993
rect 19978 59984 19984 59996
rect 20036 59984 20042 60036
rect 35161 60027 35219 60033
rect 35161 59993 35173 60027
rect 35207 60024 35219 60027
rect 35802 60024 35808 60036
rect 35207 59996 35808 60024
rect 35207 59993 35219 59996
rect 35161 59987 35219 59993
rect 35802 59984 35808 59996
rect 35860 59984 35866 60036
rect 36262 60024 36268 60036
rect 36223 59996 36268 60024
rect 36262 59984 36268 59996
rect 36320 59984 36326 60036
rect 38120 60024 38148 60055
rect 41046 60052 41052 60064
rect 41104 60052 41110 60104
rect 56318 60052 56324 60104
rect 56376 60092 56382 60104
rect 62945 60095 63003 60101
rect 62945 60092 62957 60095
rect 56376 60064 62957 60092
rect 56376 60052 56382 60064
rect 62945 60061 62957 60064
rect 62991 60061 63003 60095
rect 62945 60055 63003 60061
rect 38930 60024 38936 60036
rect 37752 59996 38148 60024
rect 38891 59996 38936 60024
rect 37752 59968 37780 59996
rect 38930 59984 38936 59996
rect 38988 59984 38994 60036
rect 40497 60027 40555 60033
rect 40497 59993 40509 60027
rect 40543 60024 40555 60027
rect 40586 60024 40592 60036
rect 40543 59996 40592 60024
rect 40543 59993 40555 59996
rect 40497 59987 40555 59993
rect 40586 59984 40592 59996
rect 40644 59984 40650 60036
rect 77754 60024 77760 60036
rect 45526 59996 64874 60024
rect 77715 59996 77760 60024
rect 1486 59916 1492 59968
rect 1544 59956 1550 59968
rect 1949 59959 2007 59965
rect 1949 59956 1961 59959
rect 1544 59928 1961 59956
rect 1544 59916 1550 59928
rect 1949 59925 1961 59928
rect 1995 59925 2007 59959
rect 1949 59919 2007 59925
rect 35253 59959 35311 59965
rect 35253 59925 35265 59959
rect 35299 59956 35311 59959
rect 35342 59956 35348 59968
rect 35299 59928 35348 59956
rect 35299 59925 35311 59928
rect 35253 59919 35311 59925
rect 35342 59916 35348 59928
rect 35400 59916 35406 59968
rect 37734 59956 37740 59968
rect 37695 59928 37740 59956
rect 37734 59916 37740 59928
rect 37792 59916 37798 59968
rect 39209 59959 39267 59965
rect 39209 59925 39221 59959
rect 39255 59956 39267 59959
rect 45526 59956 45554 59996
rect 63034 59956 63040 59968
rect 39255 59928 45554 59956
rect 62995 59928 63040 59956
rect 39255 59925 39267 59928
rect 39209 59919 39267 59925
rect 63034 59916 63040 59928
rect 63092 59916 63098 59968
rect 64846 59956 64874 59996
rect 77754 59984 77760 59996
rect 77812 59984 77818 60036
rect 77478 59956 77484 59968
rect 64846 59928 77484 59956
rect 77478 59916 77484 59928
rect 77536 59916 77542 59968
rect 1104 59866 78844 59888
rect 1104 59814 19574 59866
rect 19626 59814 19638 59866
rect 19690 59814 19702 59866
rect 19754 59814 19766 59866
rect 19818 59814 19830 59866
rect 19882 59814 50294 59866
rect 50346 59814 50358 59866
rect 50410 59814 50422 59866
rect 50474 59814 50486 59866
rect 50538 59814 50550 59866
rect 50602 59814 78844 59866
rect 1104 59792 78844 59814
rect 4614 59712 4620 59764
rect 4672 59752 4678 59764
rect 4672 59724 26234 59752
rect 4672 59712 4678 59724
rect 26206 59684 26234 59724
rect 33134 59712 33140 59764
rect 33192 59752 33198 59764
rect 36262 59752 36268 59764
rect 33192 59724 36268 59752
rect 33192 59712 33198 59724
rect 36262 59712 36268 59724
rect 36320 59712 36326 59764
rect 77754 59752 77760 59764
rect 77715 59724 77760 59752
rect 77754 59712 77760 59724
rect 77812 59712 77818 59764
rect 37734 59684 37740 59696
rect 26206 59656 37740 59684
rect 37734 59644 37740 59656
rect 37792 59644 37798 59696
rect 1946 59576 1952 59628
rect 2004 59616 2010 59628
rect 38657 59619 38715 59625
rect 38657 59616 38669 59619
rect 2004 59588 38669 59616
rect 2004 59576 2010 59588
rect 38657 59585 38669 59588
rect 38703 59616 38715 59619
rect 38933 59619 38991 59625
rect 38933 59616 38945 59619
rect 38703 59588 38945 59616
rect 38703 59585 38715 59588
rect 38657 59579 38715 59585
rect 38933 59585 38945 59588
rect 38979 59585 38991 59619
rect 38933 59579 38991 59585
rect 39574 59576 39580 59628
rect 39632 59616 39638 59628
rect 39945 59619 40003 59625
rect 39945 59616 39957 59619
rect 39632 59588 39957 59616
rect 39632 59576 39638 59588
rect 39945 59585 39957 59588
rect 39991 59585 40003 59619
rect 39945 59579 40003 59585
rect 41049 59619 41107 59625
rect 41049 59585 41061 59619
rect 41095 59616 41107 59619
rect 41138 59616 41144 59628
rect 41095 59588 41144 59616
rect 41095 59585 41107 59588
rect 41049 59579 41107 59585
rect 41138 59576 41144 59588
rect 41196 59576 41202 59628
rect 71314 59576 71320 59628
rect 71372 59616 71378 59628
rect 74721 59619 74779 59625
rect 74721 59616 74733 59619
rect 71372 59588 74733 59616
rect 71372 59576 71378 59588
rect 74721 59585 74733 59588
rect 74767 59585 74779 59619
rect 77938 59616 77944 59628
rect 77899 59588 77944 59616
rect 74721 59579 74779 59585
rect 77938 59576 77944 59588
rect 77996 59576 78002 59628
rect 39114 59548 39120 59560
rect 39075 59520 39120 59548
rect 39114 59508 39120 59520
rect 39172 59508 39178 59560
rect 40497 59551 40555 59557
rect 40497 59517 40509 59551
rect 40543 59548 40555 59551
rect 77386 59548 77392 59560
rect 40543 59520 77392 59548
rect 40543 59517 40555 59520
rect 40497 59511 40555 59517
rect 77386 59508 77392 59520
rect 77444 59508 77450 59560
rect 41233 59483 41291 59489
rect 41233 59480 41245 59483
rect 26206 59452 41245 59480
rect 1394 59372 1400 59424
rect 1452 59412 1458 59424
rect 26206 59412 26234 59452
rect 41233 59449 41245 59452
rect 41279 59449 41291 59483
rect 41233 59443 41291 59449
rect 1452 59384 26234 59412
rect 74537 59415 74595 59421
rect 1452 59372 1458 59384
rect 74537 59381 74549 59415
rect 74583 59412 74595 59415
rect 77386 59412 77392 59424
rect 74583 59384 77392 59412
rect 74583 59381 74595 59384
rect 74537 59375 74595 59381
rect 77386 59372 77392 59384
rect 77444 59372 77450 59424
rect 1104 59322 78844 59344
rect 1104 59270 4214 59322
rect 4266 59270 4278 59322
rect 4330 59270 4342 59322
rect 4394 59270 4406 59322
rect 4458 59270 4470 59322
rect 4522 59270 34934 59322
rect 34986 59270 34998 59322
rect 35050 59270 35062 59322
rect 35114 59270 35126 59322
rect 35178 59270 35190 59322
rect 35242 59270 65654 59322
rect 65706 59270 65718 59322
rect 65770 59270 65782 59322
rect 65834 59270 65846 59322
rect 65898 59270 65910 59322
rect 65962 59270 78844 59322
rect 1104 59248 78844 59270
rect 2958 59208 2964 59220
rect 2919 59180 2964 59208
rect 2958 59168 2964 59180
rect 3016 59168 3022 59220
rect 1394 59004 1400 59016
rect 1355 58976 1400 59004
rect 1394 58964 1400 58976
rect 1452 58964 1458 59016
rect 2777 59007 2835 59013
rect 2777 58973 2789 59007
rect 2823 59004 2835 59007
rect 2958 59004 2964 59016
rect 2823 58976 2964 59004
rect 2823 58973 2835 58976
rect 2777 58967 2835 58973
rect 2958 58964 2964 58976
rect 3016 58964 3022 59016
rect 39666 58964 39672 59016
rect 39724 59004 39730 59016
rect 39853 59007 39911 59013
rect 39853 59004 39865 59007
rect 39724 58976 39865 59004
rect 39724 58964 39730 58976
rect 39853 58973 39865 58976
rect 39899 58973 39911 59007
rect 39853 58967 39911 58973
rect 40129 58939 40187 58945
rect 40129 58905 40141 58939
rect 40175 58936 40187 58939
rect 63862 58936 63868 58948
rect 40175 58908 63868 58936
rect 40175 58905 40187 58908
rect 40129 58899 40187 58905
rect 63862 58896 63868 58908
rect 63920 58896 63926 58948
rect 1578 58868 1584 58880
rect 1539 58840 1584 58868
rect 1578 58828 1584 58840
rect 1636 58828 1642 58880
rect 1104 58778 78844 58800
rect 1104 58726 19574 58778
rect 19626 58726 19638 58778
rect 19690 58726 19702 58778
rect 19754 58726 19766 58778
rect 19818 58726 19830 58778
rect 19882 58726 50294 58778
rect 50346 58726 50358 58778
rect 50410 58726 50422 58778
rect 50474 58726 50486 58778
rect 50538 58726 50550 58778
rect 50602 58726 78844 58778
rect 1104 58704 78844 58726
rect 1394 58624 1400 58676
rect 1452 58664 1458 58676
rect 2777 58667 2835 58673
rect 2777 58664 2789 58667
rect 1452 58636 2789 58664
rect 1452 58624 1458 58636
rect 2777 58633 2789 58636
rect 2823 58633 2835 58667
rect 2777 58627 2835 58633
rect 1670 58488 1676 58540
rect 1728 58488 1734 58540
rect 2958 58528 2964 58540
rect 2919 58500 2964 58528
rect 2958 58488 2964 58500
rect 3016 58488 3022 58540
rect 1688 58336 1716 58488
rect 1670 58284 1676 58336
rect 1728 58284 1734 58336
rect 1104 58234 78844 58256
rect 1104 58182 4214 58234
rect 4266 58182 4278 58234
rect 4330 58182 4342 58234
rect 4394 58182 4406 58234
rect 4458 58182 4470 58234
rect 4522 58182 34934 58234
rect 34986 58182 34998 58234
rect 35050 58182 35062 58234
rect 35114 58182 35126 58234
rect 35178 58182 35190 58234
rect 35242 58182 65654 58234
rect 65706 58182 65718 58234
rect 65770 58182 65782 58234
rect 65834 58182 65846 58234
rect 65898 58182 65910 58234
rect 65962 58182 78844 58234
rect 1104 58160 78844 58182
rect 1104 57690 78844 57712
rect 1104 57638 19574 57690
rect 19626 57638 19638 57690
rect 19690 57638 19702 57690
rect 19754 57638 19766 57690
rect 19818 57638 19830 57690
rect 19882 57638 50294 57690
rect 50346 57638 50358 57690
rect 50410 57638 50422 57690
rect 50474 57638 50486 57690
rect 50538 57638 50550 57690
rect 50602 57638 78844 57690
rect 1104 57616 78844 57638
rect 1104 57146 78844 57168
rect 1104 57094 4214 57146
rect 4266 57094 4278 57146
rect 4330 57094 4342 57146
rect 4394 57094 4406 57146
rect 4458 57094 4470 57146
rect 4522 57094 34934 57146
rect 34986 57094 34998 57146
rect 35050 57094 35062 57146
rect 35114 57094 35126 57146
rect 35178 57094 35190 57146
rect 35242 57094 65654 57146
rect 65706 57094 65718 57146
rect 65770 57094 65782 57146
rect 65834 57094 65846 57146
rect 65898 57094 65910 57146
rect 65962 57094 78844 57146
rect 1104 57072 78844 57094
rect 1104 56602 78844 56624
rect 1104 56550 19574 56602
rect 19626 56550 19638 56602
rect 19690 56550 19702 56602
rect 19754 56550 19766 56602
rect 19818 56550 19830 56602
rect 19882 56550 50294 56602
rect 50346 56550 50358 56602
rect 50410 56550 50422 56602
rect 50474 56550 50486 56602
rect 50538 56550 50550 56602
rect 50602 56550 78844 56602
rect 1104 56528 78844 56550
rect 77665 56355 77723 56361
rect 77665 56321 77677 56355
rect 77711 56352 77723 56355
rect 77754 56352 77760 56364
rect 77711 56324 77760 56352
rect 77711 56321 77723 56324
rect 77665 56315 77723 56321
rect 77754 56312 77760 56324
rect 77812 56312 77818 56364
rect 77846 56148 77852 56160
rect 77807 56120 77852 56148
rect 77846 56108 77852 56120
rect 77904 56108 77910 56160
rect 1104 56058 78844 56080
rect 1104 56006 4214 56058
rect 4266 56006 4278 56058
rect 4330 56006 4342 56058
rect 4394 56006 4406 56058
rect 4458 56006 4470 56058
rect 4522 56006 34934 56058
rect 34986 56006 34998 56058
rect 35050 56006 35062 56058
rect 35114 56006 35126 56058
rect 35178 56006 35190 56058
rect 35242 56006 65654 56058
rect 65706 56006 65718 56058
rect 65770 56006 65782 56058
rect 65834 56006 65846 56058
rect 65898 56006 65910 56058
rect 65962 56006 78844 56058
rect 1104 55984 78844 56006
rect 1104 55514 78844 55536
rect 1104 55462 19574 55514
rect 19626 55462 19638 55514
rect 19690 55462 19702 55514
rect 19754 55462 19766 55514
rect 19818 55462 19830 55514
rect 19882 55462 50294 55514
rect 50346 55462 50358 55514
rect 50410 55462 50422 55514
rect 50474 55462 50486 55514
rect 50538 55462 50550 55514
rect 50602 55462 78844 55514
rect 1104 55440 78844 55462
rect 1104 54970 78844 54992
rect 1104 54918 4214 54970
rect 4266 54918 4278 54970
rect 4330 54918 4342 54970
rect 4394 54918 4406 54970
rect 4458 54918 4470 54970
rect 4522 54918 34934 54970
rect 34986 54918 34998 54970
rect 35050 54918 35062 54970
rect 35114 54918 35126 54970
rect 35178 54918 35190 54970
rect 35242 54918 65654 54970
rect 65706 54918 65718 54970
rect 65770 54918 65782 54970
rect 65834 54918 65846 54970
rect 65898 54918 65910 54970
rect 65962 54918 78844 54970
rect 1104 54896 78844 54918
rect 1673 54655 1731 54661
rect 1673 54621 1685 54655
rect 1719 54652 1731 54655
rect 2041 54655 2099 54661
rect 2041 54652 2053 54655
rect 1719 54624 2053 54652
rect 1719 54621 1731 54624
rect 1673 54615 1731 54621
rect 2041 54621 2053 54624
rect 2087 54652 2099 54655
rect 40494 54652 40500 54664
rect 2087 54624 40500 54652
rect 2087 54621 2099 54624
rect 2041 54615 2099 54621
rect 40494 54612 40500 54624
rect 40552 54612 40558 54664
rect 1486 54516 1492 54528
rect 1447 54488 1492 54516
rect 1486 54476 1492 54488
rect 1544 54476 1550 54528
rect 1104 54426 78844 54448
rect 1104 54374 19574 54426
rect 19626 54374 19638 54426
rect 19690 54374 19702 54426
rect 19754 54374 19766 54426
rect 19818 54374 19830 54426
rect 19882 54374 50294 54426
rect 50346 54374 50358 54426
rect 50410 54374 50422 54426
rect 50474 54374 50486 54426
rect 50538 54374 50550 54426
rect 50602 54374 78844 54426
rect 1104 54352 78844 54374
rect 1104 53882 78844 53904
rect 1104 53830 4214 53882
rect 4266 53830 4278 53882
rect 4330 53830 4342 53882
rect 4394 53830 4406 53882
rect 4458 53830 4470 53882
rect 4522 53830 34934 53882
rect 34986 53830 34998 53882
rect 35050 53830 35062 53882
rect 35114 53830 35126 53882
rect 35178 53830 35190 53882
rect 35242 53830 65654 53882
rect 65706 53830 65718 53882
rect 65770 53830 65782 53882
rect 65834 53830 65846 53882
rect 65898 53830 65910 53882
rect 65962 53830 78844 53882
rect 1104 53808 78844 53830
rect 1104 53338 78844 53360
rect 1104 53286 19574 53338
rect 19626 53286 19638 53338
rect 19690 53286 19702 53338
rect 19754 53286 19766 53338
rect 19818 53286 19830 53338
rect 19882 53286 50294 53338
rect 50346 53286 50358 53338
rect 50410 53286 50422 53338
rect 50474 53286 50486 53338
rect 50538 53286 50550 53338
rect 50602 53286 78844 53338
rect 1104 53264 78844 53286
rect 1104 52794 78844 52816
rect 1104 52742 4214 52794
rect 4266 52742 4278 52794
rect 4330 52742 4342 52794
rect 4394 52742 4406 52794
rect 4458 52742 4470 52794
rect 4522 52742 34934 52794
rect 34986 52742 34998 52794
rect 35050 52742 35062 52794
rect 35114 52742 35126 52794
rect 35178 52742 35190 52794
rect 35242 52742 65654 52794
rect 65706 52742 65718 52794
rect 65770 52742 65782 52794
rect 65834 52742 65846 52794
rect 65898 52742 65910 52794
rect 65962 52742 78844 52794
rect 1104 52720 78844 52742
rect 1104 52250 78844 52272
rect 1104 52198 19574 52250
rect 19626 52198 19638 52250
rect 19690 52198 19702 52250
rect 19754 52198 19766 52250
rect 19818 52198 19830 52250
rect 19882 52198 50294 52250
rect 50346 52198 50358 52250
rect 50410 52198 50422 52250
rect 50474 52198 50486 52250
rect 50538 52198 50550 52250
rect 50602 52198 78844 52250
rect 1104 52176 78844 52198
rect 77386 51960 77392 52012
rect 77444 52000 77450 52012
rect 77665 52003 77723 52009
rect 77665 52000 77677 52003
rect 77444 51972 77677 52000
rect 77444 51960 77450 51972
rect 77665 51969 77677 51972
rect 77711 51969 77723 52003
rect 77665 51963 77723 51969
rect 77846 51796 77852 51808
rect 77807 51768 77852 51796
rect 77846 51756 77852 51768
rect 77904 51756 77910 51808
rect 1104 51706 78844 51728
rect 1104 51654 4214 51706
rect 4266 51654 4278 51706
rect 4330 51654 4342 51706
rect 4394 51654 4406 51706
rect 4458 51654 4470 51706
rect 4522 51654 34934 51706
rect 34986 51654 34998 51706
rect 35050 51654 35062 51706
rect 35114 51654 35126 51706
rect 35178 51654 35190 51706
rect 35242 51654 65654 51706
rect 65706 51654 65718 51706
rect 65770 51654 65782 51706
rect 65834 51654 65846 51706
rect 65898 51654 65910 51706
rect 65962 51654 78844 51706
rect 1104 51632 78844 51654
rect 1104 51162 78844 51184
rect 1104 51110 19574 51162
rect 19626 51110 19638 51162
rect 19690 51110 19702 51162
rect 19754 51110 19766 51162
rect 19818 51110 19830 51162
rect 19882 51110 50294 51162
rect 50346 51110 50358 51162
rect 50410 51110 50422 51162
rect 50474 51110 50486 51162
rect 50538 51110 50550 51162
rect 50602 51110 78844 51162
rect 1104 51088 78844 51110
rect 1673 50915 1731 50921
rect 1673 50881 1685 50915
rect 1719 50912 1731 50915
rect 2041 50915 2099 50921
rect 2041 50912 2053 50915
rect 1719 50884 2053 50912
rect 1719 50881 1731 50884
rect 1673 50875 1731 50881
rect 2041 50881 2053 50884
rect 2087 50912 2099 50915
rect 39482 50912 39488 50924
rect 2087 50884 39488 50912
rect 2087 50881 2099 50884
rect 2041 50875 2099 50881
rect 39482 50872 39488 50884
rect 39540 50872 39546 50924
rect 1486 50708 1492 50720
rect 1447 50680 1492 50708
rect 1486 50668 1492 50680
rect 1544 50668 1550 50720
rect 1104 50618 78844 50640
rect 1104 50566 4214 50618
rect 4266 50566 4278 50618
rect 4330 50566 4342 50618
rect 4394 50566 4406 50618
rect 4458 50566 4470 50618
rect 4522 50566 34934 50618
rect 34986 50566 34998 50618
rect 35050 50566 35062 50618
rect 35114 50566 35126 50618
rect 35178 50566 35190 50618
rect 35242 50566 65654 50618
rect 65706 50566 65718 50618
rect 65770 50566 65782 50618
rect 65834 50566 65846 50618
rect 65898 50566 65910 50618
rect 65962 50566 78844 50618
rect 1104 50544 78844 50566
rect 1104 50074 78844 50096
rect 1104 50022 19574 50074
rect 19626 50022 19638 50074
rect 19690 50022 19702 50074
rect 19754 50022 19766 50074
rect 19818 50022 19830 50074
rect 19882 50022 50294 50074
rect 50346 50022 50358 50074
rect 50410 50022 50422 50074
rect 50474 50022 50486 50074
rect 50538 50022 50550 50074
rect 50602 50022 78844 50074
rect 1104 50000 78844 50022
rect 1104 49530 78844 49552
rect 1104 49478 4214 49530
rect 4266 49478 4278 49530
rect 4330 49478 4342 49530
rect 4394 49478 4406 49530
rect 4458 49478 4470 49530
rect 4522 49478 34934 49530
rect 34986 49478 34998 49530
rect 35050 49478 35062 49530
rect 35114 49478 35126 49530
rect 35178 49478 35190 49530
rect 35242 49478 65654 49530
rect 65706 49478 65718 49530
rect 65770 49478 65782 49530
rect 65834 49478 65846 49530
rect 65898 49478 65910 49530
rect 65962 49478 78844 49530
rect 1104 49456 78844 49478
rect 1104 48986 78844 49008
rect 1104 48934 19574 48986
rect 19626 48934 19638 48986
rect 19690 48934 19702 48986
rect 19754 48934 19766 48986
rect 19818 48934 19830 48986
rect 19882 48934 50294 48986
rect 50346 48934 50358 48986
rect 50410 48934 50422 48986
rect 50474 48934 50486 48986
rect 50538 48934 50550 48986
rect 50602 48934 78844 48986
rect 1104 48912 78844 48934
rect 1104 48442 78844 48464
rect 1104 48390 4214 48442
rect 4266 48390 4278 48442
rect 4330 48390 4342 48442
rect 4394 48390 4406 48442
rect 4458 48390 4470 48442
rect 4522 48390 34934 48442
rect 34986 48390 34998 48442
rect 35050 48390 35062 48442
rect 35114 48390 35126 48442
rect 35178 48390 35190 48442
rect 35242 48390 65654 48442
rect 65706 48390 65718 48442
rect 65770 48390 65782 48442
rect 65834 48390 65846 48442
rect 65898 48390 65910 48442
rect 65962 48390 78844 48442
rect 1104 48368 78844 48390
rect 39850 48220 39856 48272
rect 39908 48260 39914 48272
rect 75822 48260 75828 48272
rect 39908 48232 75828 48260
rect 39908 48220 39914 48232
rect 75822 48220 75828 48232
rect 75880 48220 75886 48272
rect 1104 47898 78844 47920
rect 1104 47846 19574 47898
rect 19626 47846 19638 47898
rect 19690 47846 19702 47898
rect 19754 47846 19766 47898
rect 19818 47846 19830 47898
rect 19882 47846 50294 47898
rect 50346 47846 50358 47898
rect 50410 47846 50422 47898
rect 50474 47846 50486 47898
rect 50538 47846 50550 47898
rect 50602 47846 78844 47898
rect 1104 47824 78844 47846
rect 1104 47354 78844 47376
rect 1104 47302 4214 47354
rect 4266 47302 4278 47354
rect 4330 47302 4342 47354
rect 4394 47302 4406 47354
rect 4458 47302 4470 47354
rect 4522 47302 34934 47354
rect 34986 47302 34998 47354
rect 35050 47302 35062 47354
rect 35114 47302 35126 47354
rect 35178 47302 35190 47354
rect 35242 47302 65654 47354
rect 65706 47302 65718 47354
rect 65770 47302 65782 47354
rect 65834 47302 65846 47354
rect 65898 47302 65910 47354
rect 65962 47302 78844 47354
rect 1104 47280 78844 47302
rect 1578 47172 1584 47184
rect 1539 47144 1584 47172
rect 1578 47132 1584 47144
rect 1636 47132 1642 47184
rect 1397 47039 1455 47045
rect 1397 47005 1409 47039
rect 1443 47036 1455 47039
rect 2866 47036 2872 47048
rect 1443 47008 2872 47036
rect 1443 47005 1455 47008
rect 1397 46999 1455 47005
rect 2866 46996 2872 47008
rect 2924 46996 2930 47048
rect 1104 46810 78844 46832
rect 1104 46758 19574 46810
rect 19626 46758 19638 46810
rect 19690 46758 19702 46810
rect 19754 46758 19766 46810
rect 19818 46758 19830 46810
rect 19882 46758 50294 46810
rect 50346 46758 50358 46810
rect 50410 46758 50422 46810
rect 50474 46758 50486 46810
rect 50538 46758 50550 46810
rect 50602 46758 78844 46810
rect 1104 46736 78844 46758
rect 1104 46266 78844 46288
rect 1104 46214 4214 46266
rect 4266 46214 4278 46266
rect 4330 46214 4342 46266
rect 4394 46214 4406 46266
rect 4458 46214 4470 46266
rect 4522 46214 34934 46266
rect 34986 46214 34998 46266
rect 35050 46214 35062 46266
rect 35114 46214 35126 46266
rect 35178 46214 35190 46266
rect 35242 46214 65654 46266
rect 65706 46214 65718 46266
rect 65770 46214 65782 46266
rect 65834 46214 65846 46266
rect 65898 46214 65910 46266
rect 65962 46214 78844 46266
rect 1104 46192 78844 46214
rect 1104 45722 78844 45744
rect 1104 45670 19574 45722
rect 19626 45670 19638 45722
rect 19690 45670 19702 45722
rect 19754 45670 19766 45722
rect 19818 45670 19830 45722
rect 19882 45670 50294 45722
rect 50346 45670 50358 45722
rect 50410 45670 50422 45722
rect 50474 45670 50486 45722
rect 50538 45670 50550 45722
rect 50602 45670 78844 45722
rect 1104 45648 78844 45670
rect 1104 45178 78844 45200
rect 1104 45126 4214 45178
rect 4266 45126 4278 45178
rect 4330 45126 4342 45178
rect 4394 45126 4406 45178
rect 4458 45126 4470 45178
rect 4522 45126 34934 45178
rect 34986 45126 34998 45178
rect 35050 45126 35062 45178
rect 35114 45126 35126 45178
rect 35178 45126 35190 45178
rect 35242 45126 65654 45178
rect 65706 45126 65718 45178
rect 65770 45126 65782 45178
rect 65834 45126 65846 45178
rect 65898 45126 65910 45178
rect 65962 45126 78844 45178
rect 1104 45104 78844 45126
rect 1104 44634 78844 44656
rect 1104 44582 19574 44634
rect 19626 44582 19638 44634
rect 19690 44582 19702 44634
rect 19754 44582 19766 44634
rect 19818 44582 19830 44634
rect 19882 44582 50294 44634
rect 50346 44582 50358 44634
rect 50410 44582 50422 44634
rect 50474 44582 50486 44634
rect 50538 44582 50550 44634
rect 50602 44582 78844 44634
rect 1104 44560 78844 44582
rect 1104 44090 78844 44112
rect 1104 44038 4214 44090
rect 4266 44038 4278 44090
rect 4330 44038 4342 44090
rect 4394 44038 4406 44090
rect 4458 44038 4470 44090
rect 4522 44038 34934 44090
rect 34986 44038 34998 44090
rect 35050 44038 35062 44090
rect 35114 44038 35126 44090
rect 35178 44038 35190 44090
rect 35242 44038 65654 44090
rect 65706 44038 65718 44090
rect 65770 44038 65782 44090
rect 65834 44038 65846 44090
rect 65898 44038 65910 44090
rect 65962 44038 78844 44090
rect 1104 44016 78844 44038
rect 76558 43732 76564 43784
rect 76616 43772 76622 43784
rect 77849 43775 77907 43781
rect 77849 43772 77861 43775
rect 76616 43744 77861 43772
rect 76616 43732 76622 43744
rect 77849 43741 77861 43744
rect 77895 43741 77907 43775
rect 77849 43735 77907 43741
rect 78030 43636 78036 43648
rect 77991 43608 78036 43636
rect 78030 43596 78036 43608
rect 78088 43596 78094 43648
rect 1104 43546 78844 43568
rect 1104 43494 19574 43546
rect 19626 43494 19638 43546
rect 19690 43494 19702 43546
rect 19754 43494 19766 43546
rect 19818 43494 19830 43546
rect 19882 43494 50294 43546
rect 50346 43494 50358 43546
rect 50410 43494 50422 43546
rect 50474 43494 50486 43546
rect 50538 43494 50550 43546
rect 50602 43494 78844 43546
rect 1104 43472 78844 43494
rect 1854 43296 1860 43308
rect 1815 43268 1860 43296
rect 1854 43256 1860 43268
rect 1912 43256 1918 43308
rect 2133 43095 2191 43101
rect 2133 43061 2145 43095
rect 2179 43092 2191 43095
rect 39574 43092 39580 43104
rect 2179 43064 39580 43092
rect 2179 43061 2191 43064
rect 2133 43055 2191 43061
rect 39574 43052 39580 43064
rect 39632 43052 39638 43104
rect 1104 43002 78844 43024
rect 1104 42950 4214 43002
rect 4266 42950 4278 43002
rect 4330 42950 4342 43002
rect 4394 42950 4406 43002
rect 4458 42950 4470 43002
rect 4522 42950 34934 43002
rect 34986 42950 34998 43002
rect 35050 42950 35062 43002
rect 35114 42950 35126 43002
rect 35178 42950 35190 43002
rect 35242 42950 65654 43002
rect 65706 42950 65718 43002
rect 65770 42950 65782 43002
rect 65834 42950 65846 43002
rect 65898 42950 65910 43002
rect 65962 42950 78844 43002
rect 1104 42928 78844 42950
rect 77754 42752 77760 42764
rect 77715 42724 77760 42752
rect 77754 42712 77760 42724
rect 77812 42712 77818 42764
rect 77570 42616 77576 42628
rect 77531 42588 77576 42616
rect 77570 42576 77576 42588
rect 77628 42576 77634 42628
rect 1104 42458 78844 42480
rect 1104 42406 19574 42458
rect 19626 42406 19638 42458
rect 19690 42406 19702 42458
rect 19754 42406 19766 42458
rect 19818 42406 19830 42458
rect 19882 42406 50294 42458
rect 50346 42406 50358 42458
rect 50410 42406 50422 42458
rect 50474 42406 50486 42458
rect 50538 42406 50550 42458
rect 50602 42406 78844 42458
rect 1104 42384 78844 42406
rect 1104 41914 78844 41936
rect 1104 41862 4214 41914
rect 4266 41862 4278 41914
rect 4330 41862 4342 41914
rect 4394 41862 4406 41914
rect 4458 41862 4470 41914
rect 4522 41862 34934 41914
rect 34986 41862 34998 41914
rect 35050 41862 35062 41914
rect 35114 41862 35126 41914
rect 35178 41862 35190 41914
rect 35242 41862 65654 41914
rect 65706 41862 65718 41914
rect 65770 41862 65782 41914
rect 65834 41862 65846 41914
rect 65898 41862 65910 41914
rect 65962 41862 78844 41914
rect 1104 41840 78844 41862
rect 1104 41370 78844 41392
rect 1104 41318 19574 41370
rect 19626 41318 19638 41370
rect 19690 41318 19702 41370
rect 19754 41318 19766 41370
rect 19818 41318 19830 41370
rect 19882 41318 50294 41370
rect 50346 41318 50358 41370
rect 50410 41318 50422 41370
rect 50474 41318 50486 41370
rect 50538 41318 50550 41370
rect 50602 41318 78844 41370
rect 1104 41296 78844 41318
rect 1104 40826 78844 40848
rect 1104 40774 4214 40826
rect 4266 40774 4278 40826
rect 4330 40774 4342 40826
rect 4394 40774 4406 40826
rect 4458 40774 4470 40826
rect 4522 40774 34934 40826
rect 34986 40774 34998 40826
rect 35050 40774 35062 40826
rect 35114 40774 35126 40826
rect 35178 40774 35190 40826
rect 35242 40774 65654 40826
rect 65706 40774 65718 40826
rect 65770 40774 65782 40826
rect 65834 40774 65846 40826
rect 65898 40774 65910 40826
rect 65962 40774 78844 40826
rect 1104 40752 78844 40774
rect 77478 40468 77484 40520
rect 77536 40508 77542 40520
rect 77849 40511 77907 40517
rect 77849 40508 77861 40511
rect 77536 40480 77861 40508
rect 77536 40468 77542 40480
rect 77849 40477 77861 40480
rect 77895 40477 77907 40511
rect 77849 40471 77907 40477
rect 78030 40372 78036 40384
rect 77991 40344 78036 40372
rect 78030 40332 78036 40344
rect 78088 40332 78094 40384
rect 1104 40282 78844 40304
rect 1104 40230 19574 40282
rect 19626 40230 19638 40282
rect 19690 40230 19702 40282
rect 19754 40230 19766 40282
rect 19818 40230 19830 40282
rect 19882 40230 50294 40282
rect 50346 40230 50358 40282
rect 50410 40230 50422 40282
rect 50474 40230 50486 40282
rect 50538 40230 50550 40282
rect 50602 40230 78844 40282
rect 1104 40208 78844 40230
rect 77478 40168 77484 40180
rect 77439 40140 77484 40168
rect 77478 40128 77484 40140
rect 77536 40128 77542 40180
rect 77570 40060 77576 40112
rect 77628 40100 77634 40112
rect 77628 40072 77708 40100
rect 77628 40060 77634 40072
rect 77680 40041 77708 40072
rect 77665 40035 77723 40041
rect 77665 40001 77677 40035
rect 77711 40001 77723 40035
rect 77665 39995 77723 40001
rect 1104 39738 78844 39760
rect 1104 39686 4214 39738
rect 4266 39686 4278 39738
rect 4330 39686 4342 39738
rect 4394 39686 4406 39738
rect 4458 39686 4470 39738
rect 4522 39686 34934 39738
rect 34986 39686 34998 39738
rect 35050 39686 35062 39738
rect 35114 39686 35126 39738
rect 35178 39686 35190 39738
rect 35242 39686 65654 39738
rect 65706 39686 65718 39738
rect 65770 39686 65782 39738
rect 65834 39686 65846 39738
rect 65898 39686 65910 39738
rect 65962 39686 78844 39738
rect 1104 39664 78844 39686
rect 1104 39194 78844 39216
rect 1104 39142 19574 39194
rect 19626 39142 19638 39194
rect 19690 39142 19702 39194
rect 19754 39142 19766 39194
rect 19818 39142 19830 39194
rect 19882 39142 50294 39194
rect 50346 39142 50358 39194
rect 50410 39142 50422 39194
rect 50474 39142 50486 39194
rect 50538 39142 50550 39194
rect 50602 39142 78844 39194
rect 1104 39120 78844 39142
rect 1854 38944 1860 38956
rect 1815 38916 1860 38944
rect 1854 38904 1860 38916
rect 1912 38904 1918 38956
rect 2133 38743 2191 38749
rect 2133 38709 2145 38743
rect 2179 38740 2191 38743
rect 38838 38740 38844 38752
rect 2179 38712 38844 38740
rect 2179 38709 2191 38712
rect 2133 38703 2191 38709
rect 38838 38700 38844 38712
rect 38896 38700 38902 38752
rect 1104 38650 78844 38672
rect 1104 38598 4214 38650
rect 4266 38598 4278 38650
rect 4330 38598 4342 38650
rect 4394 38598 4406 38650
rect 4458 38598 4470 38650
rect 4522 38598 34934 38650
rect 34986 38598 34998 38650
rect 35050 38598 35062 38650
rect 35114 38598 35126 38650
rect 35178 38598 35190 38650
rect 35242 38598 65654 38650
rect 65706 38598 65718 38650
rect 65770 38598 65782 38650
rect 65834 38598 65846 38650
rect 65898 38598 65910 38650
rect 65962 38598 78844 38650
rect 1104 38576 78844 38598
rect 1104 38106 78844 38128
rect 1104 38054 19574 38106
rect 19626 38054 19638 38106
rect 19690 38054 19702 38106
rect 19754 38054 19766 38106
rect 19818 38054 19830 38106
rect 19882 38054 50294 38106
rect 50346 38054 50358 38106
rect 50410 38054 50422 38106
rect 50474 38054 50486 38106
rect 50538 38054 50550 38106
rect 50602 38054 78844 38106
rect 1104 38032 78844 38054
rect 1104 37562 78844 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 34934 37562
rect 34986 37510 34998 37562
rect 35050 37510 35062 37562
rect 35114 37510 35126 37562
rect 35178 37510 35190 37562
rect 35242 37510 65654 37562
rect 65706 37510 65718 37562
rect 65770 37510 65782 37562
rect 65834 37510 65846 37562
rect 65898 37510 65910 37562
rect 65962 37510 78844 37562
rect 1104 37488 78844 37510
rect 1104 37018 78844 37040
rect 1104 36966 19574 37018
rect 19626 36966 19638 37018
rect 19690 36966 19702 37018
rect 19754 36966 19766 37018
rect 19818 36966 19830 37018
rect 19882 36966 50294 37018
rect 50346 36966 50358 37018
rect 50410 36966 50422 37018
rect 50474 36966 50486 37018
rect 50538 36966 50550 37018
rect 50602 36966 78844 37018
rect 1104 36944 78844 36966
rect 1104 36474 78844 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 65654 36474
rect 65706 36422 65718 36474
rect 65770 36422 65782 36474
rect 65834 36422 65846 36474
rect 65898 36422 65910 36474
rect 65962 36422 78844 36474
rect 1104 36400 78844 36422
rect 77846 36156 77852 36168
rect 77807 36128 77852 36156
rect 77846 36116 77852 36128
rect 77904 36116 77910 36168
rect 78030 36020 78036 36032
rect 77991 35992 78036 36020
rect 78030 35980 78036 35992
rect 78088 35980 78094 36032
rect 1104 35930 78844 35952
rect 1104 35878 19574 35930
rect 19626 35878 19638 35930
rect 19690 35878 19702 35930
rect 19754 35878 19766 35930
rect 19818 35878 19830 35930
rect 19882 35878 50294 35930
rect 50346 35878 50358 35930
rect 50410 35878 50422 35930
rect 50474 35878 50486 35930
rect 50538 35878 50550 35930
rect 50602 35878 78844 35930
rect 1104 35856 78844 35878
rect 1104 35386 78844 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 65654 35386
rect 65706 35334 65718 35386
rect 65770 35334 65782 35386
rect 65834 35334 65846 35386
rect 65898 35334 65910 35386
rect 65962 35334 78844 35386
rect 1104 35312 78844 35334
rect 1397 35071 1455 35077
rect 1397 35037 1409 35071
rect 1443 35068 1455 35071
rect 1486 35068 1492 35080
rect 1443 35040 1492 35068
rect 1443 35037 1455 35040
rect 1397 35031 1455 35037
rect 1486 35028 1492 35040
rect 1544 35028 1550 35080
rect 1578 34932 1584 34944
rect 1539 34904 1584 34932
rect 1578 34892 1584 34904
rect 1636 34892 1642 34944
rect 1104 34842 78844 34864
rect 1104 34790 19574 34842
rect 19626 34790 19638 34842
rect 19690 34790 19702 34842
rect 19754 34790 19766 34842
rect 19818 34790 19830 34842
rect 19882 34790 50294 34842
rect 50346 34790 50358 34842
rect 50410 34790 50422 34842
rect 50474 34790 50486 34842
rect 50538 34790 50550 34842
rect 50602 34790 78844 34842
rect 1104 34768 78844 34790
rect 71869 34663 71927 34669
rect 71869 34629 71881 34663
rect 71915 34660 71927 34663
rect 76558 34660 76564 34672
rect 71915 34632 76564 34660
rect 71915 34629 71927 34632
rect 71869 34623 71927 34629
rect 76558 34620 76564 34632
rect 76616 34620 76622 34672
rect 66622 34552 66628 34604
rect 66680 34592 66686 34604
rect 71685 34595 71743 34601
rect 71685 34592 71697 34595
rect 66680 34564 71697 34592
rect 66680 34552 66686 34564
rect 71685 34561 71697 34564
rect 71731 34561 71743 34595
rect 71685 34555 71743 34561
rect 1104 34298 78844 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 65654 34298
rect 65706 34246 65718 34298
rect 65770 34246 65782 34298
rect 65834 34246 65846 34298
rect 65898 34246 65910 34298
rect 65962 34246 78844 34298
rect 1104 34224 78844 34246
rect 1104 33754 78844 33776
rect 1104 33702 19574 33754
rect 19626 33702 19638 33754
rect 19690 33702 19702 33754
rect 19754 33702 19766 33754
rect 19818 33702 19830 33754
rect 19882 33702 50294 33754
rect 50346 33702 50358 33754
rect 50410 33702 50422 33754
rect 50474 33702 50486 33754
rect 50538 33702 50550 33754
rect 50602 33702 78844 33754
rect 1104 33680 78844 33702
rect 1104 33210 78844 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 65654 33210
rect 65706 33158 65718 33210
rect 65770 33158 65782 33210
rect 65834 33158 65846 33210
rect 65898 33158 65910 33210
rect 65962 33158 78844 33210
rect 1104 33136 78844 33158
rect 77846 33096 77852 33108
rect 77807 33068 77852 33096
rect 77846 33056 77852 33068
rect 77904 33056 77910 33108
rect 78030 32892 78036 32904
rect 77991 32864 78036 32892
rect 78030 32852 78036 32864
rect 78088 32852 78094 32904
rect 1104 32666 78844 32688
rect 1104 32614 19574 32666
rect 19626 32614 19638 32666
rect 19690 32614 19702 32666
rect 19754 32614 19766 32666
rect 19818 32614 19830 32666
rect 19882 32614 50294 32666
rect 50346 32614 50358 32666
rect 50410 32614 50422 32666
rect 50474 32614 50486 32666
rect 50538 32614 50550 32666
rect 50602 32614 78844 32666
rect 1104 32592 78844 32614
rect 77665 32419 77723 32425
rect 77665 32385 77677 32419
rect 77711 32416 77723 32419
rect 77754 32416 77760 32428
rect 77711 32388 77760 32416
rect 77711 32385 77723 32388
rect 77665 32379 77723 32385
rect 77754 32376 77760 32388
rect 77812 32376 77818 32428
rect 77846 32212 77852 32224
rect 77807 32184 77852 32212
rect 77846 32172 77852 32184
rect 77904 32172 77910 32224
rect 1104 32122 78844 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 65654 32122
rect 65706 32070 65718 32122
rect 65770 32070 65782 32122
rect 65834 32070 65846 32122
rect 65898 32070 65910 32122
rect 65962 32070 78844 32122
rect 1104 32048 78844 32070
rect 1673 31875 1731 31881
rect 1673 31841 1685 31875
rect 1719 31872 1731 31875
rect 40770 31872 40776 31884
rect 1719 31844 40776 31872
rect 1719 31841 1731 31844
rect 1673 31835 1731 31841
rect 40770 31832 40776 31844
rect 40828 31832 40834 31884
rect 1394 31804 1400 31816
rect 1355 31776 1400 31804
rect 1394 31764 1400 31776
rect 1452 31764 1458 31816
rect 1104 31578 78844 31600
rect 1104 31526 19574 31578
rect 19626 31526 19638 31578
rect 19690 31526 19702 31578
rect 19754 31526 19766 31578
rect 19818 31526 19830 31578
rect 19882 31526 50294 31578
rect 50346 31526 50358 31578
rect 50410 31526 50422 31578
rect 50474 31526 50486 31578
rect 50538 31526 50550 31578
rect 50602 31526 78844 31578
rect 1104 31504 78844 31526
rect 1104 31034 78844 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 65654 31034
rect 65706 30982 65718 31034
rect 65770 30982 65782 31034
rect 65834 30982 65846 31034
rect 65898 30982 65910 31034
rect 65962 30982 78844 31034
rect 1104 30960 78844 30982
rect 1104 30490 78844 30512
rect 1104 30438 19574 30490
rect 19626 30438 19638 30490
rect 19690 30438 19702 30490
rect 19754 30438 19766 30490
rect 19818 30438 19830 30490
rect 19882 30438 50294 30490
rect 50346 30438 50358 30490
rect 50410 30438 50422 30490
rect 50474 30438 50486 30490
rect 50538 30438 50550 30490
rect 50602 30438 78844 30490
rect 1104 30416 78844 30438
rect 1104 29946 78844 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 65654 29946
rect 65706 29894 65718 29946
rect 65770 29894 65782 29946
rect 65834 29894 65846 29946
rect 65898 29894 65910 29946
rect 65962 29894 78844 29946
rect 1104 29872 78844 29894
rect 1104 29402 78844 29424
rect 1104 29350 19574 29402
rect 19626 29350 19638 29402
rect 19690 29350 19702 29402
rect 19754 29350 19766 29402
rect 19818 29350 19830 29402
rect 19882 29350 50294 29402
rect 50346 29350 50358 29402
rect 50410 29350 50422 29402
rect 50474 29350 50486 29402
rect 50538 29350 50550 29402
rect 50602 29350 78844 29402
rect 1104 29328 78844 29350
rect 1104 28858 78844 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 65654 28858
rect 65706 28806 65718 28858
rect 65770 28806 65782 28858
rect 65834 28806 65846 28858
rect 65898 28806 65910 28858
rect 65962 28806 78844 28858
rect 1104 28784 78844 28806
rect 1104 28314 78844 28336
rect 1104 28262 19574 28314
rect 19626 28262 19638 28314
rect 19690 28262 19702 28314
rect 19754 28262 19766 28314
rect 19818 28262 19830 28314
rect 19882 28262 50294 28314
rect 50346 28262 50358 28314
rect 50410 28262 50422 28314
rect 50474 28262 50486 28314
rect 50538 28262 50550 28314
rect 50602 28262 78844 28314
rect 1104 28240 78844 28262
rect 77757 28203 77815 28209
rect 77757 28169 77769 28203
rect 77803 28200 77815 28203
rect 78030 28200 78036 28212
rect 77803 28172 78036 28200
rect 77803 28169 77815 28172
rect 77757 28163 77815 28169
rect 78030 28160 78036 28172
rect 78088 28160 78094 28212
rect 77938 28064 77944 28076
rect 77899 28036 77944 28064
rect 77938 28024 77944 28036
rect 77996 28024 78002 28076
rect 1104 27770 78844 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 65654 27770
rect 65706 27718 65718 27770
rect 65770 27718 65782 27770
rect 65834 27718 65846 27770
rect 65898 27718 65910 27770
rect 65962 27718 78844 27770
rect 1104 27696 78844 27718
rect 1394 27452 1400 27464
rect 1355 27424 1400 27452
rect 1394 27412 1400 27424
rect 1452 27412 1458 27464
rect 1673 27387 1731 27393
rect 1673 27353 1685 27387
rect 1719 27384 1731 27387
rect 39666 27384 39672 27396
rect 1719 27356 39672 27384
rect 1719 27353 1731 27356
rect 1673 27347 1731 27353
rect 39666 27344 39672 27356
rect 39724 27344 39730 27396
rect 1104 27226 78844 27248
rect 1104 27174 19574 27226
rect 19626 27174 19638 27226
rect 19690 27174 19702 27226
rect 19754 27174 19766 27226
rect 19818 27174 19830 27226
rect 19882 27174 50294 27226
rect 50346 27174 50358 27226
rect 50410 27174 50422 27226
rect 50474 27174 50486 27226
rect 50538 27174 50550 27226
rect 50602 27174 78844 27226
rect 1104 27152 78844 27174
rect 1104 26682 78844 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 65654 26682
rect 65706 26630 65718 26682
rect 65770 26630 65782 26682
rect 65834 26630 65846 26682
rect 65898 26630 65910 26682
rect 65962 26630 78844 26682
rect 1104 26608 78844 26630
rect 1104 26138 78844 26160
rect 1104 26086 19574 26138
rect 19626 26086 19638 26138
rect 19690 26086 19702 26138
rect 19754 26086 19766 26138
rect 19818 26086 19830 26138
rect 19882 26086 50294 26138
rect 50346 26086 50358 26138
rect 50410 26086 50422 26138
rect 50474 26086 50486 26138
rect 50538 26086 50550 26138
rect 50602 26086 78844 26138
rect 1104 26064 78844 26086
rect 39577 25891 39635 25897
rect 39577 25857 39589 25891
rect 39623 25888 39635 25891
rect 40221 25891 40279 25897
rect 40221 25888 40233 25891
rect 39623 25860 40233 25888
rect 39623 25857 39635 25860
rect 39577 25851 39635 25857
rect 40221 25857 40233 25860
rect 40267 25888 40279 25891
rect 77846 25888 77852 25900
rect 40267 25860 77852 25888
rect 40267 25857 40279 25860
rect 40221 25851 40279 25857
rect 77846 25848 77852 25860
rect 77904 25848 77910 25900
rect 39574 25644 39580 25696
rect 39632 25684 39638 25696
rect 39945 25687 40003 25693
rect 39945 25684 39957 25687
rect 39632 25656 39957 25684
rect 39632 25644 39638 25656
rect 39945 25653 39957 25656
rect 39991 25653 40003 25687
rect 39945 25647 40003 25653
rect 1104 25594 78844 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 65654 25594
rect 65706 25542 65718 25594
rect 65770 25542 65782 25594
rect 65834 25542 65846 25594
rect 65898 25542 65910 25594
rect 65962 25542 78844 25594
rect 1104 25520 78844 25542
rect 1762 25440 1768 25492
rect 1820 25480 1826 25492
rect 39574 25480 39580 25492
rect 1820 25452 39580 25480
rect 1820 25440 1826 25452
rect 39574 25440 39580 25452
rect 39632 25440 39638 25492
rect 1104 25050 78844 25072
rect 1104 24998 19574 25050
rect 19626 24998 19638 25050
rect 19690 24998 19702 25050
rect 19754 24998 19766 25050
rect 19818 24998 19830 25050
rect 19882 24998 50294 25050
rect 50346 24998 50358 25050
rect 50410 24998 50422 25050
rect 50474 24998 50486 25050
rect 50538 24998 50550 25050
rect 50602 24998 78844 25050
rect 1104 24976 78844 24998
rect 77665 24803 77723 24809
rect 77665 24800 77677 24803
rect 77312 24772 77677 24800
rect 39114 24556 39120 24608
rect 39172 24596 39178 24608
rect 77312 24605 77340 24772
rect 77665 24769 77677 24772
rect 77711 24769 77723 24803
rect 77665 24763 77723 24769
rect 77297 24599 77355 24605
rect 77297 24596 77309 24599
rect 39172 24568 77309 24596
rect 39172 24556 39178 24568
rect 77297 24565 77309 24568
rect 77343 24565 77355 24599
rect 77846 24596 77852 24608
rect 77807 24568 77852 24596
rect 77297 24559 77355 24565
rect 77846 24556 77852 24568
rect 77904 24556 77910 24608
rect 1104 24506 78844 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 65654 24506
rect 65706 24454 65718 24506
rect 65770 24454 65782 24506
rect 65834 24454 65846 24506
rect 65898 24454 65910 24506
rect 65962 24454 78844 24506
rect 1104 24432 78844 24454
rect 1104 23962 78844 23984
rect 1104 23910 19574 23962
rect 19626 23910 19638 23962
rect 19690 23910 19702 23962
rect 19754 23910 19766 23962
rect 19818 23910 19830 23962
rect 19882 23910 50294 23962
rect 50346 23910 50358 23962
rect 50410 23910 50422 23962
rect 50474 23910 50486 23962
rect 50538 23910 50550 23962
rect 50602 23910 78844 23962
rect 1104 23888 78844 23910
rect 1394 23712 1400 23724
rect 1355 23684 1400 23712
rect 1394 23672 1400 23684
rect 1452 23672 1458 23724
rect 1673 23647 1731 23653
rect 1673 23613 1685 23647
rect 1719 23644 1731 23647
rect 38930 23644 38936 23656
rect 1719 23616 38936 23644
rect 1719 23613 1731 23616
rect 1673 23607 1731 23613
rect 38930 23604 38936 23616
rect 38988 23604 38994 23656
rect 1104 23418 78844 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 65654 23418
rect 65706 23366 65718 23418
rect 65770 23366 65782 23418
rect 65834 23366 65846 23418
rect 65898 23366 65910 23418
rect 65962 23366 78844 23418
rect 1104 23344 78844 23366
rect 1104 22874 78844 22896
rect 1104 22822 19574 22874
rect 19626 22822 19638 22874
rect 19690 22822 19702 22874
rect 19754 22822 19766 22874
rect 19818 22822 19830 22874
rect 19882 22822 50294 22874
rect 50346 22822 50358 22874
rect 50410 22822 50422 22874
rect 50474 22822 50486 22874
rect 50538 22822 50550 22874
rect 50602 22822 78844 22874
rect 1104 22800 78844 22822
rect 1104 22330 78844 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 65654 22330
rect 65706 22278 65718 22330
rect 65770 22278 65782 22330
rect 65834 22278 65846 22330
rect 65898 22278 65910 22330
rect 65962 22278 78844 22330
rect 1104 22256 78844 22278
rect 1104 21786 78844 21808
rect 1104 21734 19574 21786
rect 19626 21734 19638 21786
rect 19690 21734 19702 21786
rect 19754 21734 19766 21786
rect 19818 21734 19830 21786
rect 19882 21734 50294 21786
rect 50346 21734 50358 21786
rect 50410 21734 50422 21786
rect 50474 21734 50486 21786
rect 50538 21734 50550 21786
rect 50602 21734 78844 21786
rect 1104 21712 78844 21734
rect 1104 21242 78844 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 65654 21242
rect 65706 21190 65718 21242
rect 65770 21190 65782 21242
rect 65834 21190 65846 21242
rect 65898 21190 65910 21242
rect 65962 21190 78844 21242
rect 1104 21168 78844 21190
rect 77754 20884 77760 20936
rect 77812 20924 77818 20936
rect 77849 20927 77907 20933
rect 77849 20924 77861 20927
rect 77812 20896 77861 20924
rect 77812 20884 77818 20896
rect 77849 20893 77861 20896
rect 77895 20893 77907 20927
rect 77849 20887 77907 20893
rect 78030 20788 78036 20800
rect 77991 20760 78036 20788
rect 78030 20748 78036 20760
rect 78088 20748 78094 20800
rect 1104 20698 78844 20720
rect 1104 20646 19574 20698
rect 19626 20646 19638 20698
rect 19690 20646 19702 20698
rect 19754 20646 19766 20698
rect 19818 20646 19830 20698
rect 19882 20646 50294 20698
rect 50346 20646 50358 20698
rect 50410 20646 50422 20698
rect 50474 20646 50486 20698
rect 50538 20646 50550 20698
rect 50602 20646 78844 20698
rect 1104 20624 78844 20646
rect 1104 20154 78844 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 65654 20154
rect 65706 20102 65718 20154
rect 65770 20102 65782 20154
rect 65834 20102 65846 20154
rect 65898 20102 65910 20154
rect 65962 20102 78844 20154
rect 1104 20080 78844 20102
rect 1104 19610 78844 19632
rect 1104 19558 19574 19610
rect 19626 19558 19638 19610
rect 19690 19558 19702 19610
rect 19754 19558 19766 19610
rect 19818 19558 19830 19610
rect 19882 19558 50294 19610
rect 50346 19558 50358 19610
rect 50410 19558 50422 19610
rect 50474 19558 50486 19610
rect 50538 19558 50550 19610
rect 50602 19558 78844 19610
rect 1104 19536 78844 19558
rect 1397 19363 1455 19369
rect 1397 19329 1409 19363
rect 1443 19360 1455 19363
rect 1486 19360 1492 19372
rect 1443 19332 1492 19360
rect 1443 19329 1455 19332
rect 1397 19323 1455 19329
rect 1486 19320 1492 19332
rect 1544 19320 1550 19372
rect 1578 19156 1584 19168
rect 1539 19128 1584 19156
rect 1578 19116 1584 19128
rect 1636 19116 1642 19168
rect 1104 19066 78844 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 65654 19066
rect 65706 19014 65718 19066
rect 65770 19014 65782 19066
rect 65834 19014 65846 19066
rect 65898 19014 65910 19066
rect 65962 19014 78844 19066
rect 1104 18992 78844 19014
rect 1104 18522 78844 18544
rect 1104 18470 19574 18522
rect 19626 18470 19638 18522
rect 19690 18470 19702 18522
rect 19754 18470 19766 18522
rect 19818 18470 19830 18522
rect 19882 18470 50294 18522
rect 50346 18470 50358 18522
rect 50410 18470 50422 18522
rect 50474 18470 50486 18522
rect 50538 18470 50550 18522
rect 50602 18470 78844 18522
rect 1104 18448 78844 18470
rect 1104 17978 78844 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 65654 17978
rect 65706 17926 65718 17978
rect 65770 17926 65782 17978
rect 65834 17926 65846 17978
rect 65898 17926 65910 17978
rect 65962 17926 78844 17978
rect 1104 17904 78844 17926
rect 1104 17434 78844 17456
rect 1104 17382 19574 17434
rect 19626 17382 19638 17434
rect 19690 17382 19702 17434
rect 19754 17382 19766 17434
rect 19818 17382 19830 17434
rect 19882 17382 50294 17434
rect 50346 17382 50358 17434
rect 50410 17382 50422 17434
rect 50474 17382 50486 17434
rect 50538 17382 50550 17434
rect 50602 17382 78844 17434
rect 1104 17360 78844 17382
rect 1104 16890 78844 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 65654 16890
rect 65706 16838 65718 16890
rect 65770 16838 65782 16890
rect 65834 16838 65846 16890
rect 65898 16838 65910 16890
rect 65962 16838 78844 16890
rect 1104 16816 78844 16838
rect 63034 16532 63040 16584
rect 63092 16572 63098 16584
rect 77849 16575 77907 16581
rect 77849 16572 77861 16575
rect 63092 16544 77861 16572
rect 63092 16532 63098 16544
rect 77849 16541 77861 16544
rect 77895 16541 77907 16575
rect 77849 16535 77907 16541
rect 78030 16436 78036 16448
rect 77991 16408 78036 16436
rect 78030 16396 78036 16408
rect 78088 16396 78094 16448
rect 1104 16346 78844 16368
rect 1104 16294 19574 16346
rect 19626 16294 19638 16346
rect 19690 16294 19702 16346
rect 19754 16294 19766 16346
rect 19818 16294 19830 16346
rect 19882 16294 50294 16346
rect 50346 16294 50358 16346
rect 50410 16294 50422 16346
rect 50474 16294 50486 16346
rect 50538 16294 50550 16346
rect 50602 16294 78844 16346
rect 1104 16272 78844 16294
rect 1762 16192 1768 16244
rect 1820 16232 1826 16244
rect 1949 16235 2007 16241
rect 1949 16232 1961 16235
rect 1820 16204 1961 16232
rect 1820 16192 1826 16204
rect 1949 16201 1961 16204
rect 1995 16201 2007 16235
rect 1949 16195 2007 16201
rect 1673 16099 1731 16105
rect 1673 16065 1685 16099
rect 1719 16096 1731 16099
rect 1780 16096 1808 16192
rect 1719 16068 1808 16096
rect 1719 16065 1731 16068
rect 1673 16059 1731 16065
rect 1486 15892 1492 15904
rect 1447 15864 1492 15892
rect 1486 15852 1492 15864
rect 1544 15852 1550 15904
rect 1104 15802 78844 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 65654 15802
rect 65706 15750 65718 15802
rect 65770 15750 65782 15802
rect 65834 15750 65846 15802
rect 65898 15750 65910 15802
rect 65962 15750 78844 15802
rect 1104 15728 78844 15750
rect 1104 15258 78844 15280
rect 1104 15206 19574 15258
rect 19626 15206 19638 15258
rect 19690 15206 19702 15258
rect 19754 15206 19766 15258
rect 19818 15206 19830 15258
rect 19882 15206 50294 15258
rect 50346 15206 50358 15258
rect 50410 15206 50422 15258
rect 50474 15206 50486 15258
rect 50538 15206 50550 15258
rect 50602 15206 78844 15258
rect 1104 15184 78844 15206
rect 1104 14714 78844 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 65654 14714
rect 65706 14662 65718 14714
rect 65770 14662 65782 14714
rect 65834 14662 65846 14714
rect 65898 14662 65910 14714
rect 65962 14662 78844 14714
rect 1104 14640 78844 14662
rect 1104 14170 78844 14192
rect 1104 14118 19574 14170
rect 19626 14118 19638 14170
rect 19690 14118 19702 14170
rect 19754 14118 19766 14170
rect 19818 14118 19830 14170
rect 19882 14118 50294 14170
rect 50346 14118 50358 14170
rect 50410 14118 50422 14170
rect 50474 14118 50486 14170
rect 50538 14118 50550 14170
rect 50602 14118 78844 14170
rect 1104 14096 78844 14118
rect 1104 13626 78844 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 65654 13626
rect 65706 13574 65718 13626
rect 65770 13574 65782 13626
rect 65834 13574 65846 13626
rect 65898 13574 65910 13626
rect 65962 13574 78844 13626
rect 1104 13552 78844 13574
rect 2866 13512 2872 13524
rect 2827 13484 2872 13512
rect 2866 13472 2872 13484
rect 2924 13472 2930 13524
rect 2406 13268 2412 13320
rect 2464 13308 2470 13320
rect 2685 13311 2743 13317
rect 2685 13308 2697 13311
rect 2464 13280 2697 13308
rect 2464 13268 2470 13280
rect 2685 13277 2697 13280
rect 2731 13277 2743 13311
rect 2685 13271 2743 13277
rect 1104 13082 78844 13104
rect 1104 13030 19574 13082
rect 19626 13030 19638 13082
rect 19690 13030 19702 13082
rect 19754 13030 19766 13082
rect 19818 13030 19830 13082
rect 19882 13030 50294 13082
rect 50346 13030 50358 13082
rect 50410 13030 50422 13082
rect 50474 13030 50486 13082
rect 50538 13030 50550 13082
rect 50602 13030 78844 13082
rect 1104 13008 78844 13030
rect 77662 12860 77668 12912
rect 77720 12900 77726 12912
rect 77757 12903 77815 12909
rect 77757 12900 77769 12903
rect 77720 12872 77769 12900
rect 77720 12860 77726 12872
rect 77757 12869 77769 12872
rect 77803 12869 77815 12903
rect 77757 12863 77815 12869
rect 77202 12792 77208 12844
rect 77260 12832 77266 12844
rect 77481 12835 77539 12841
rect 77481 12832 77493 12835
rect 77260 12804 77493 12832
rect 77260 12792 77266 12804
rect 77481 12801 77493 12804
rect 77527 12801 77539 12835
rect 77481 12795 77539 12801
rect 1104 12538 78844 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 65654 12538
rect 65706 12486 65718 12538
rect 65770 12486 65782 12538
rect 65834 12486 65846 12538
rect 65898 12486 65910 12538
rect 65962 12486 78844 12538
rect 1104 12464 78844 12486
rect 18322 12112 18328 12164
rect 18380 12152 18386 12164
rect 40313 12155 40371 12161
rect 40313 12152 40325 12155
rect 18380 12124 40325 12152
rect 18380 12112 18386 12124
rect 40313 12121 40325 12124
rect 40359 12121 40371 12155
rect 40313 12115 40371 12121
rect 40589 12087 40647 12093
rect 40589 12053 40601 12087
rect 40635 12084 40647 12087
rect 77754 12084 77760 12096
rect 40635 12056 77760 12084
rect 40635 12053 40647 12056
rect 40589 12047 40647 12053
rect 77754 12044 77760 12056
rect 77812 12044 77818 12096
rect 1104 11994 78844 12016
rect 1104 11942 19574 11994
rect 19626 11942 19638 11994
rect 19690 11942 19702 11994
rect 19754 11942 19766 11994
rect 19818 11942 19830 11994
rect 19882 11942 50294 11994
rect 50346 11942 50358 11994
rect 50410 11942 50422 11994
rect 50474 11942 50486 11994
rect 50538 11942 50550 11994
rect 50602 11942 78844 11994
rect 1104 11920 78844 11942
rect 1673 11815 1731 11821
rect 1673 11781 1685 11815
rect 1719 11812 1731 11815
rect 3050 11812 3056 11824
rect 1719 11784 3056 11812
rect 1719 11781 1731 11784
rect 1673 11775 1731 11781
rect 3050 11772 3056 11784
rect 3108 11772 3114 11824
rect 1394 11744 1400 11756
rect 1355 11716 1400 11744
rect 1394 11704 1400 11716
rect 1452 11704 1458 11756
rect 1104 11450 78844 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 65654 11450
rect 65706 11398 65718 11450
rect 65770 11398 65782 11450
rect 65834 11398 65846 11450
rect 65898 11398 65910 11450
rect 65962 11398 78844 11450
rect 1104 11376 78844 11398
rect 1104 10906 78844 10928
rect 1104 10854 19574 10906
rect 19626 10854 19638 10906
rect 19690 10854 19702 10906
rect 19754 10854 19766 10906
rect 19818 10854 19830 10906
rect 19882 10854 50294 10906
rect 50346 10854 50358 10906
rect 50410 10854 50422 10906
rect 50474 10854 50486 10906
rect 50538 10854 50550 10906
rect 50602 10854 78844 10906
rect 1104 10832 78844 10854
rect 1104 10362 78844 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 65654 10362
rect 65706 10310 65718 10362
rect 65770 10310 65782 10362
rect 65834 10310 65846 10362
rect 65898 10310 65910 10362
rect 65962 10310 78844 10362
rect 1104 10288 78844 10310
rect 78033 10115 78091 10121
rect 78033 10081 78045 10115
rect 78079 10112 78091 10115
rect 78122 10112 78128 10124
rect 78079 10084 78128 10112
rect 78079 10081 78091 10084
rect 78033 10075 78091 10081
rect 78122 10072 78128 10084
rect 78180 10072 78186 10124
rect 77481 10047 77539 10053
rect 77481 10013 77493 10047
rect 77527 10044 77539 10047
rect 77938 10044 77944 10056
rect 77527 10016 77944 10044
rect 77527 10013 77539 10016
rect 77481 10007 77539 10013
rect 77938 10004 77944 10016
rect 77996 10004 78002 10056
rect 1104 9818 78844 9840
rect 1104 9766 19574 9818
rect 19626 9766 19638 9818
rect 19690 9766 19702 9818
rect 19754 9766 19766 9818
rect 19818 9766 19830 9818
rect 19882 9766 50294 9818
rect 50346 9766 50358 9818
rect 50410 9766 50422 9818
rect 50474 9766 50486 9818
rect 50538 9766 50550 9818
rect 50602 9766 78844 9818
rect 1104 9744 78844 9766
rect 1104 9274 78844 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 65654 9274
rect 65706 9222 65718 9274
rect 65770 9222 65782 9274
rect 65834 9222 65846 9274
rect 65898 9222 65910 9274
rect 65962 9222 78844 9274
rect 1104 9200 78844 9222
rect 77849 8959 77907 8965
rect 77849 8956 77861 8959
rect 77496 8928 77861 8956
rect 40586 8780 40592 8832
rect 40644 8820 40650 8832
rect 77496 8829 77524 8928
rect 77849 8925 77861 8928
rect 77895 8925 77907 8959
rect 77849 8919 77907 8925
rect 77481 8823 77539 8829
rect 77481 8820 77493 8823
rect 40644 8792 77493 8820
rect 40644 8780 40650 8792
rect 77481 8789 77493 8792
rect 77527 8789 77539 8823
rect 78030 8820 78036 8832
rect 77991 8792 78036 8820
rect 77481 8783 77539 8789
rect 78030 8780 78036 8792
rect 78088 8780 78094 8832
rect 1104 8730 78844 8752
rect 1104 8678 19574 8730
rect 19626 8678 19638 8730
rect 19690 8678 19702 8730
rect 19754 8678 19766 8730
rect 19818 8678 19830 8730
rect 19882 8678 50294 8730
rect 50346 8678 50358 8730
rect 50410 8678 50422 8730
rect 50474 8678 50486 8730
rect 50538 8678 50550 8730
rect 50602 8678 78844 8730
rect 1104 8656 78844 8678
rect 1104 8186 78844 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 65654 8186
rect 65706 8134 65718 8186
rect 65770 8134 65782 8186
rect 65834 8134 65846 8186
rect 65898 8134 65910 8186
rect 65962 8134 78844 8186
rect 1104 8112 78844 8134
rect 1397 7871 1455 7877
rect 1397 7837 1409 7871
rect 1443 7868 1455 7871
rect 2682 7868 2688 7880
rect 1443 7840 2688 7868
rect 1443 7837 1455 7840
rect 1397 7831 1455 7837
rect 2682 7828 2688 7840
rect 2740 7828 2746 7880
rect 1578 7732 1584 7744
rect 1539 7704 1584 7732
rect 1578 7692 1584 7704
rect 1636 7692 1642 7744
rect 1104 7642 78844 7664
rect 1104 7590 19574 7642
rect 19626 7590 19638 7642
rect 19690 7590 19702 7642
rect 19754 7590 19766 7642
rect 19818 7590 19830 7642
rect 19882 7590 50294 7642
rect 50346 7590 50358 7642
rect 50410 7590 50422 7642
rect 50474 7590 50486 7642
rect 50538 7590 50550 7642
rect 50602 7590 78844 7642
rect 1104 7568 78844 7590
rect 2406 7528 2412 7540
rect 2367 7500 2412 7528
rect 2406 7488 2412 7500
rect 2464 7488 2470 7540
rect 2682 7528 2688 7540
rect 2643 7500 2688 7528
rect 2682 7488 2688 7500
rect 2740 7488 2746 7540
rect 2424 7392 2452 7488
rect 2869 7395 2927 7401
rect 2869 7392 2881 7395
rect 2424 7364 2881 7392
rect 2869 7361 2881 7364
rect 2915 7392 2927 7395
rect 29914 7392 29920 7404
rect 2915 7364 29920 7392
rect 2915 7361 2927 7364
rect 2869 7355 2927 7361
rect 29914 7352 29920 7364
rect 29972 7352 29978 7404
rect 1104 7098 78844 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 65654 7098
rect 65706 7046 65718 7098
rect 65770 7046 65782 7098
rect 65834 7046 65846 7098
rect 65898 7046 65910 7098
rect 65962 7046 78844 7098
rect 1104 7024 78844 7046
rect 1104 6554 78844 6576
rect 1104 6502 19574 6554
rect 19626 6502 19638 6554
rect 19690 6502 19702 6554
rect 19754 6502 19766 6554
rect 19818 6502 19830 6554
rect 19882 6502 50294 6554
rect 50346 6502 50358 6554
rect 50410 6502 50422 6554
rect 50474 6502 50486 6554
rect 50538 6502 50550 6554
rect 50602 6502 78844 6554
rect 1104 6480 78844 6502
rect 1104 6010 78844 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 65654 6010
rect 65706 5958 65718 6010
rect 65770 5958 65782 6010
rect 65834 5958 65846 6010
rect 65898 5958 65910 6010
rect 65962 5958 78844 6010
rect 1104 5936 78844 5958
rect 1104 5466 78844 5488
rect 1104 5414 19574 5466
rect 19626 5414 19638 5466
rect 19690 5414 19702 5466
rect 19754 5414 19766 5466
rect 19818 5414 19830 5466
rect 19882 5414 50294 5466
rect 50346 5414 50358 5466
rect 50410 5414 50422 5466
rect 50474 5414 50486 5466
rect 50538 5414 50550 5466
rect 50602 5414 78844 5466
rect 1104 5392 78844 5414
rect 77662 5216 77668 5228
rect 77623 5188 77668 5216
rect 77662 5176 77668 5188
rect 77720 5176 77726 5228
rect 77846 5012 77852 5024
rect 77807 4984 77852 5012
rect 77846 4972 77852 4984
rect 77904 4972 77910 5024
rect 1104 4922 78844 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 65654 4922
rect 65706 4870 65718 4922
rect 65770 4870 65782 4922
rect 65834 4870 65846 4922
rect 65898 4870 65910 4922
rect 65962 4870 78844 4922
rect 1104 4848 78844 4870
rect 77662 4768 77668 4820
rect 77720 4808 77726 4820
rect 77849 4811 77907 4817
rect 77849 4808 77861 4811
rect 77720 4780 77861 4808
rect 77720 4768 77726 4780
rect 77849 4777 77861 4780
rect 77895 4777 77907 4811
rect 77849 4771 77907 4777
rect 78030 4604 78036 4616
rect 77991 4576 78036 4604
rect 78030 4564 78036 4576
rect 78088 4564 78094 4616
rect 1104 4378 78844 4400
rect 1104 4326 19574 4378
rect 19626 4326 19638 4378
rect 19690 4326 19702 4378
rect 19754 4326 19766 4378
rect 19818 4326 19830 4378
rect 19882 4326 50294 4378
rect 50346 4326 50358 4378
rect 50410 4326 50422 4378
rect 50474 4326 50486 4378
rect 50538 4326 50550 4378
rect 50602 4326 78844 4378
rect 1104 4304 78844 4326
rect 1104 3834 78844 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 65654 3834
rect 65706 3782 65718 3834
rect 65770 3782 65782 3834
rect 65834 3782 65846 3834
rect 65898 3782 65910 3834
rect 65962 3782 78844 3834
rect 1104 3760 78844 3782
rect 1670 3584 1676 3596
rect 1631 3556 1676 3584
rect 1670 3544 1676 3556
rect 1728 3544 1734 3596
rect 1394 3516 1400 3528
rect 1355 3488 1400 3516
rect 1394 3476 1400 3488
rect 1452 3476 1458 3528
rect 12434 3476 12440 3528
rect 12492 3516 12498 3528
rect 15105 3519 15163 3525
rect 15105 3516 15117 3519
rect 12492 3488 15117 3516
rect 12492 3476 12498 3488
rect 15105 3485 15117 3488
rect 15151 3485 15163 3519
rect 40954 3516 40960 3528
rect 40915 3488 40960 3516
rect 15105 3479 15163 3485
rect 40954 3476 40960 3488
rect 41012 3476 41018 3528
rect 41877 3519 41935 3525
rect 41877 3485 41889 3519
rect 41923 3516 41935 3519
rect 43898 3516 43904 3528
rect 41923 3488 43904 3516
rect 41923 3485 41935 3488
rect 41877 3479 41935 3485
rect 43898 3476 43904 3488
rect 43956 3476 43962 3528
rect 40313 3451 40371 3457
rect 40313 3417 40325 3451
rect 40359 3448 40371 3451
rect 57974 3448 57980 3460
rect 40359 3420 57980 3448
rect 40359 3417 40371 3420
rect 40313 3411 40371 3417
rect 57974 3408 57980 3420
rect 58032 3408 58038 3460
rect 14921 3383 14979 3389
rect 14921 3349 14933 3383
rect 14967 3380 14979 3383
rect 16206 3380 16212 3392
rect 14967 3352 16212 3380
rect 14967 3349 14979 3352
rect 14921 3343 14979 3349
rect 16206 3340 16212 3352
rect 16264 3340 16270 3392
rect 40402 3380 40408 3392
rect 40363 3352 40408 3380
rect 40402 3340 40408 3352
rect 40460 3340 40466 3392
rect 41138 3380 41144 3392
rect 41099 3352 41144 3380
rect 41138 3340 41144 3352
rect 41196 3340 41202 3392
rect 41690 3380 41696 3392
rect 41651 3352 41696 3380
rect 41690 3340 41696 3352
rect 41748 3340 41754 3392
rect 1104 3290 78844 3312
rect 1104 3238 19574 3290
rect 19626 3238 19638 3290
rect 19690 3238 19702 3290
rect 19754 3238 19766 3290
rect 19818 3238 19830 3290
rect 19882 3238 50294 3290
rect 50346 3238 50358 3290
rect 50410 3238 50422 3290
rect 50474 3238 50486 3290
rect 50538 3238 50550 3290
rect 50602 3238 78844 3290
rect 1104 3216 78844 3238
rect 11514 3136 11520 3188
rect 11572 3176 11578 3188
rect 40402 3176 40408 3188
rect 11572 3148 40408 3176
rect 11572 3136 11578 3148
rect 40402 3136 40408 3148
rect 40460 3136 40466 3188
rect 77297 3043 77355 3049
rect 77297 3009 77309 3043
rect 77343 3040 77355 3043
rect 77662 3040 77668 3052
rect 77343 3012 77668 3040
rect 77343 3009 77355 3012
rect 77297 3003 77355 3009
rect 77662 3000 77668 3012
rect 77720 3000 77726 3052
rect 41230 2932 41236 2984
rect 41288 2972 41294 2984
rect 77573 2975 77631 2981
rect 77573 2972 77585 2975
rect 41288 2944 77585 2972
rect 41288 2932 41294 2944
rect 77573 2941 77585 2944
rect 77619 2941 77631 2975
rect 77573 2935 77631 2941
rect 1104 2746 78844 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 65654 2746
rect 65706 2694 65718 2746
rect 65770 2694 65782 2746
rect 65834 2694 65846 2746
rect 65898 2694 65910 2746
rect 65962 2694 78844 2746
rect 1104 2672 78844 2694
rect 18322 2632 18328 2644
rect 18283 2604 18328 2632
rect 18322 2592 18328 2604
rect 18380 2592 18386 2644
rect 29914 2632 29920 2644
rect 29875 2604 29920 2632
rect 29914 2592 29920 2604
rect 29972 2592 29978 2644
rect 33134 2632 33140 2644
rect 33095 2604 33140 2632
rect 33134 2592 33140 2604
rect 33192 2592 33198 2644
rect 40954 2632 40960 2644
rect 35866 2604 40960 2632
rect 12434 2564 12440 2576
rect 1688 2536 12440 2564
rect 1688 2505 1716 2536
rect 12434 2524 12440 2536
rect 12492 2524 12498 2576
rect 15197 2567 15255 2573
rect 15197 2533 15209 2567
rect 15243 2564 15255 2567
rect 35866 2564 35894 2604
rect 40954 2592 40960 2604
rect 41012 2592 41018 2644
rect 43898 2592 43904 2644
rect 43956 2632 43962 2644
rect 47765 2635 47823 2641
rect 47765 2632 47777 2635
rect 43956 2604 47777 2632
rect 43956 2592 43962 2604
rect 47765 2601 47777 2604
rect 47811 2601 47823 2635
rect 55766 2632 55772 2644
rect 47765 2595 47823 2601
rect 50356 2604 55772 2632
rect 15243 2536 35894 2564
rect 15243 2533 15255 2536
rect 15197 2527 15255 2533
rect 41046 2524 41052 2576
rect 41104 2564 41110 2576
rect 50356 2564 50384 2604
rect 55766 2592 55772 2604
rect 55824 2592 55830 2644
rect 66622 2632 66628 2644
rect 66583 2604 66628 2632
rect 66622 2592 66628 2604
rect 66680 2592 66686 2644
rect 41104 2536 50384 2564
rect 41104 2524 41110 2536
rect 50614 2524 50620 2576
rect 50672 2564 50678 2576
rect 50672 2536 71176 2564
rect 50672 2524 50678 2536
rect 1673 2499 1731 2505
rect 1673 2465 1685 2499
rect 1719 2465 1731 2499
rect 1673 2459 1731 2465
rect 4433 2499 4491 2505
rect 4433 2465 4445 2499
rect 4479 2496 4491 2499
rect 4614 2496 4620 2508
rect 4479 2468 4620 2496
rect 4479 2465 4491 2468
rect 4433 2459 4491 2465
rect 4614 2456 4620 2468
rect 4672 2456 4678 2508
rect 19978 2456 19984 2508
rect 20036 2496 20042 2508
rect 20036 2468 25912 2496
rect 20036 2456 20042 2468
rect 14 2388 20 2440
rect 72 2428 78 2440
rect 1397 2431 1455 2437
rect 1397 2428 1409 2431
rect 72 2400 1409 2428
rect 72 2388 78 2400
rect 1397 2397 1409 2400
rect 1443 2397 1455 2431
rect 1397 2391 1455 2397
rect 3234 2388 3240 2440
rect 3292 2428 3298 2440
rect 3881 2431 3939 2437
rect 3881 2428 3893 2431
rect 3292 2400 3893 2428
rect 3292 2388 3298 2400
rect 3881 2397 3893 2400
rect 3927 2397 3939 2431
rect 3881 2391 3939 2397
rect 7098 2388 7104 2440
rect 7156 2428 7162 2440
rect 7285 2431 7343 2437
rect 7285 2428 7297 2431
rect 7156 2400 7297 2428
rect 7156 2388 7162 2400
rect 7285 2397 7297 2400
rect 7331 2397 7343 2431
rect 11514 2428 11520 2440
rect 11475 2400 11520 2428
rect 7285 2391 7343 2397
rect 11514 2388 11520 2400
rect 11572 2388 11578 2440
rect 16206 2388 16212 2440
rect 16264 2428 16270 2440
rect 25884 2437 25912 2468
rect 41138 2456 41144 2508
rect 41196 2496 41202 2508
rect 71148 2505 71176 2536
rect 71133 2499 71191 2505
rect 41196 2468 70992 2496
rect 41196 2456 41202 2468
rect 22005 2431 22063 2437
rect 22005 2428 22017 2431
rect 16264 2400 22017 2428
rect 16264 2388 16270 2400
rect 22005 2397 22017 2400
rect 22051 2397 22063 2431
rect 22005 2391 22063 2397
rect 25869 2431 25927 2437
rect 25869 2397 25881 2431
rect 25915 2397 25927 2431
rect 25869 2391 25927 2397
rect 29638 2388 29644 2440
rect 29696 2428 29702 2440
rect 29733 2431 29791 2437
rect 29733 2428 29745 2431
rect 29696 2400 29745 2428
rect 29696 2388 29702 2400
rect 29733 2397 29745 2400
rect 29779 2397 29791 2431
rect 29733 2391 29791 2397
rect 35342 2388 35348 2440
rect 35400 2428 35406 2440
rect 37277 2431 37335 2437
rect 37277 2428 37289 2431
rect 35400 2400 37289 2428
rect 35400 2388 35406 2400
rect 37277 2397 37289 2400
rect 37323 2397 37335 2431
rect 37277 2391 37335 2397
rect 40681 2431 40739 2437
rect 40681 2397 40693 2431
rect 40727 2428 40739 2431
rect 41690 2428 41696 2440
rect 40727 2400 41696 2428
rect 40727 2397 40739 2400
rect 40681 2391 40739 2397
rect 41690 2388 41696 2400
rect 41748 2388 41754 2440
rect 44450 2388 44456 2440
rect 44508 2428 44514 2440
rect 45005 2431 45063 2437
rect 45005 2428 45017 2431
rect 44508 2400 45017 2428
rect 44508 2388 44514 2400
rect 45005 2397 45017 2400
rect 45051 2397 45063 2431
rect 45005 2391 45063 2397
rect 47670 2388 47676 2440
rect 47728 2428 47734 2440
rect 47949 2431 48007 2437
rect 47949 2428 47961 2431
rect 47728 2400 47961 2428
rect 47728 2388 47734 2400
rect 47949 2397 47961 2400
rect 47995 2397 48007 2431
rect 47949 2391 48007 2397
rect 51534 2388 51540 2440
rect 51592 2428 51598 2440
rect 51629 2431 51687 2437
rect 51629 2428 51641 2431
rect 51592 2400 51641 2428
rect 51592 2388 51598 2400
rect 51629 2397 51641 2400
rect 51675 2397 51687 2431
rect 51629 2391 51687 2397
rect 55398 2388 55404 2440
rect 55456 2428 55462 2440
rect 55493 2431 55551 2437
rect 55493 2428 55505 2431
rect 55456 2400 55505 2428
rect 55456 2388 55462 2400
rect 55493 2397 55505 2400
rect 55539 2397 55551 2431
rect 55766 2428 55772 2440
rect 55727 2400 55772 2428
rect 55493 2391 55551 2397
rect 55766 2388 55772 2400
rect 55824 2388 55830 2440
rect 59081 2431 59139 2437
rect 59081 2397 59093 2431
rect 59127 2428 59139 2431
rect 59262 2428 59268 2440
rect 59127 2400 59268 2428
rect 59127 2397 59139 2400
rect 59081 2391 59139 2397
rect 59262 2388 59268 2400
rect 59320 2388 59326 2440
rect 59357 2431 59415 2437
rect 59357 2397 59369 2431
rect 59403 2397 59415 2431
rect 59357 2391 59415 2397
rect 7834 2360 7840 2372
rect 7795 2332 7840 2360
rect 7834 2320 7840 2332
rect 7892 2320 7898 2372
rect 14826 2320 14832 2372
rect 14884 2360 14890 2372
rect 15013 2363 15071 2369
rect 15013 2360 15025 2363
rect 14884 2332 15025 2360
rect 14884 2320 14890 2332
rect 15013 2329 15025 2332
rect 15059 2329 15071 2363
rect 15013 2323 15071 2329
rect 18046 2320 18052 2372
rect 18104 2360 18110 2372
rect 18233 2363 18291 2369
rect 18233 2360 18245 2363
rect 18104 2332 18245 2360
rect 18104 2320 18110 2332
rect 18233 2329 18245 2332
rect 18279 2329 18291 2363
rect 18233 2323 18291 2329
rect 32858 2320 32864 2372
rect 32916 2360 32922 2372
rect 33045 2363 33103 2369
rect 33045 2360 33057 2363
rect 32916 2332 33057 2360
rect 32916 2320 32922 2332
rect 33045 2329 33057 2332
rect 33091 2329 33103 2363
rect 33045 2323 33103 2329
rect 39758 2320 39764 2372
rect 39816 2360 39822 2372
rect 45281 2363 45339 2369
rect 45281 2360 45293 2363
rect 39816 2332 45293 2360
rect 39816 2320 39822 2332
rect 45281 2329 45293 2332
rect 45327 2329 45339 2363
rect 51902 2360 51908 2372
rect 51863 2332 51908 2360
rect 45281 2323 45339 2329
rect 51902 2320 51908 2332
rect 51960 2320 51966 2372
rect 57974 2320 57980 2372
rect 58032 2360 58038 2372
rect 59372 2360 59400 2391
rect 62482 2388 62488 2440
rect 62540 2428 62546 2440
rect 63037 2431 63095 2437
rect 63037 2428 63049 2431
rect 62540 2400 63049 2428
rect 62540 2388 62546 2400
rect 63037 2397 63049 2400
rect 63083 2397 63095 2431
rect 63037 2391 63095 2397
rect 66346 2388 66352 2440
rect 66404 2428 66410 2440
rect 66441 2431 66499 2437
rect 66441 2428 66453 2431
rect 66404 2400 66453 2428
rect 66404 2388 66410 2400
rect 66441 2397 66453 2400
rect 66487 2397 66499 2431
rect 66441 2391 66499 2397
rect 70210 2388 70216 2440
rect 70268 2428 70274 2440
rect 70857 2431 70915 2437
rect 70857 2428 70869 2431
rect 70268 2400 70869 2428
rect 70268 2388 70274 2400
rect 70857 2397 70869 2400
rect 70903 2397 70915 2431
rect 70964 2428 70992 2468
rect 71133 2465 71145 2499
rect 71179 2465 71191 2499
rect 71133 2459 71191 2465
rect 77389 2499 77447 2505
rect 77389 2465 77401 2499
rect 77435 2496 77447 2499
rect 78030 2496 78036 2508
rect 77435 2468 78036 2496
rect 77435 2465 77447 2468
rect 77389 2459 77447 2465
rect 78030 2456 78036 2468
rect 78088 2456 78094 2508
rect 73801 2431 73859 2437
rect 73801 2428 73813 2431
rect 70964 2400 73813 2428
rect 70857 2391 70915 2397
rect 73801 2397 73813 2400
rect 73847 2428 73859 2431
rect 74169 2431 74227 2437
rect 74169 2428 74181 2431
rect 73847 2400 74181 2428
rect 73847 2397 73859 2400
rect 73801 2391 73859 2397
rect 74169 2397 74181 2400
rect 74215 2397 74227 2431
rect 74169 2391 74227 2397
rect 77113 2431 77171 2437
rect 77113 2397 77125 2431
rect 77159 2428 77171 2431
rect 77294 2428 77300 2440
rect 77159 2400 77300 2428
rect 77159 2397 77171 2400
rect 77113 2391 77171 2397
rect 77294 2388 77300 2400
rect 77352 2388 77358 2440
rect 63862 2360 63868 2372
rect 58032 2332 59400 2360
rect 63823 2332 63868 2360
rect 58032 2320 58038 2332
rect 63862 2320 63868 2332
rect 63920 2320 63926 2372
rect 10962 2252 10968 2304
rect 11020 2292 11026 2304
rect 11701 2295 11759 2301
rect 11701 2292 11713 2295
rect 11020 2264 11713 2292
rect 11020 2252 11026 2264
rect 11701 2261 11713 2264
rect 11747 2261 11759 2295
rect 11701 2255 11759 2261
rect 21910 2252 21916 2304
rect 21968 2292 21974 2304
rect 22189 2295 22247 2301
rect 22189 2292 22201 2295
rect 21968 2264 22201 2292
rect 21968 2252 21974 2264
rect 22189 2261 22201 2264
rect 22235 2261 22247 2295
rect 22189 2255 22247 2261
rect 25774 2252 25780 2304
rect 25832 2292 25838 2304
rect 26053 2295 26111 2301
rect 26053 2292 26065 2295
rect 25832 2264 26065 2292
rect 25832 2252 25838 2264
rect 26053 2261 26065 2264
rect 26099 2261 26111 2295
rect 26053 2255 26111 2261
rect 36722 2252 36728 2304
rect 36780 2292 36786 2304
rect 37461 2295 37519 2301
rect 37461 2292 37473 2295
rect 36780 2264 37473 2292
rect 36780 2252 36786 2264
rect 37461 2261 37473 2264
rect 37507 2261 37519 2295
rect 37461 2255 37519 2261
rect 40586 2252 40592 2304
rect 40644 2292 40650 2304
rect 40865 2295 40923 2301
rect 40865 2292 40877 2295
rect 40644 2264 40877 2292
rect 40644 2252 40650 2264
rect 40865 2261 40877 2264
rect 40911 2261 40923 2295
rect 40865 2255 40923 2261
rect 40954 2252 40960 2304
rect 41012 2292 41018 2304
rect 50614 2292 50620 2304
rect 41012 2264 50620 2292
rect 41012 2252 41018 2264
rect 50614 2252 50620 2264
rect 50672 2252 50678 2304
rect 74074 2252 74080 2304
rect 74132 2292 74138 2304
rect 74353 2295 74411 2301
rect 74353 2292 74365 2295
rect 74132 2264 74365 2292
rect 74132 2252 74138 2264
rect 74353 2261 74365 2264
rect 74399 2261 74411 2295
rect 74353 2255 74411 2261
rect 1104 2202 78844 2224
rect 1104 2150 19574 2202
rect 19626 2150 19638 2202
rect 19690 2150 19702 2202
rect 19754 2150 19766 2202
rect 19818 2150 19830 2202
rect 19882 2150 50294 2202
rect 50346 2150 50358 2202
rect 50410 2150 50422 2202
rect 50474 2150 50486 2202
rect 50538 2150 50550 2202
rect 50602 2150 78844 2202
rect 1104 2128 78844 2150
rect 2958 1980 2964 2032
rect 3016 2020 3022 2032
rect 63862 2020 63868 2032
rect 3016 1992 63868 2020
rect 3016 1980 3022 1992
rect 63862 1980 63868 1992
rect 63920 1980 63926 2032
rect 39942 1912 39948 1964
rect 40000 1952 40006 1964
rect 51902 1952 51908 1964
rect 40000 1924 51908 1952
rect 40000 1912 40006 1924
rect 51902 1912 51908 1924
rect 51960 1912 51966 1964
rect 7834 1844 7840 1896
rect 7892 1884 7898 1896
rect 77570 1884 77576 1896
rect 7892 1856 77576 1884
rect 7892 1844 7898 1856
rect 77570 1844 77576 1856
rect 77628 1844 77634 1896
<< via1 >>
rect 19574 117478 19626 117530
rect 19638 117478 19690 117530
rect 19702 117478 19754 117530
rect 19766 117478 19818 117530
rect 19830 117478 19882 117530
rect 50294 117478 50346 117530
rect 50358 117478 50410 117530
rect 50422 117478 50474 117530
rect 50486 117478 50538 117530
rect 50550 117478 50602 117530
rect 4620 117351 4672 117360
rect 4620 117317 4629 117351
rect 4629 117317 4663 117351
rect 4663 117317 4672 117351
rect 4620 117308 4672 117317
rect 664 117240 716 117292
rect 7840 117283 7892 117292
rect 7840 117249 7849 117283
rect 7849 117249 7883 117283
rect 7883 117249 7892 117283
rect 7840 117240 7892 117249
rect 11704 117283 11756 117292
rect 11704 117249 11713 117283
rect 11713 117249 11747 117283
rect 11747 117249 11756 117283
rect 11704 117240 11756 117249
rect 15568 117283 15620 117292
rect 15568 117249 15577 117283
rect 15577 117249 15611 117283
rect 15611 117249 15620 117283
rect 15568 117240 15620 117249
rect 19432 117283 19484 117292
rect 19432 117249 19441 117283
rect 19441 117249 19475 117283
rect 19475 117249 19484 117283
rect 19432 117240 19484 117249
rect 22652 117283 22704 117292
rect 22652 117249 22661 117283
rect 22661 117249 22695 117283
rect 22695 117249 22704 117283
rect 22652 117240 22704 117249
rect 26424 117240 26476 117292
rect 28264 117240 28316 117292
rect 34704 117283 34756 117292
rect 34704 117249 34713 117283
rect 34713 117249 34747 117283
rect 34747 117249 34756 117283
rect 34704 117240 34756 117249
rect 36360 117240 36412 117292
rect 40684 117240 40736 117292
rect 45192 117283 45244 117292
rect 45192 117249 45201 117283
rect 45201 117249 45235 117283
rect 45235 117249 45244 117283
rect 45192 117240 45244 117249
rect 49240 117283 49292 117292
rect 49240 117249 49249 117283
rect 49249 117249 49283 117283
rect 49283 117249 49292 117283
rect 49240 117240 49292 117249
rect 56140 117283 56192 117292
rect 11888 117215 11940 117224
rect 11888 117181 11897 117215
rect 11897 117181 11931 117215
rect 11931 117181 11940 117215
rect 11888 117172 11940 117181
rect 35808 117172 35860 117224
rect 19340 117104 19392 117156
rect 22836 117147 22888 117156
rect 22836 117113 22845 117147
rect 22845 117113 22879 117147
rect 22879 117113 22888 117147
rect 22836 117104 22888 117113
rect 30380 117104 30432 117156
rect 34520 117104 34572 117156
rect 2320 117036 2372 117088
rect 8024 117079 8076 117088
rect 8024 117045 8033 117079
rect 8033 117045 8067 117079
rect 8067 117045 8076 117079
rect 8024 117036 8076 117045
rect 15752 117079 15804 117088
rect 15752 117045 15761 117079
rect 15761 117045 15795 117079
rect 15795 117045 15804 117079
rect 15752 117036 15804 117045
rect 37464 117104 37516 117156
rect 37648 117147 37700 117156
rect 37648 117113 37657 117147
rect 37657 117113 37691 117147
rect 37691 117113 37700 117147
rect 37648 117104 37700 117113
rect 45376 117147 45428 117156
rect 45376 117113 45385 117147
rect 45385 117113 45419 117147
rect 45419 117113 45428 117147
rect 45376 117104 45428 117113
rect 52460 117104 52512 117156
rect 56140 117249 56149 117283
rect 56149 117249 56183 117283
rect 56183 117249 56192 117283
rect 56140 117240 56192 117249
rect 59912 117240 59964 117292
rect 63868 117283 63920 117292
rect 63868 117249 63877 117283
rect 63877 117249 63911 117283
rect 63911 117249 63920 117283
rect 63868 117240 63920 117249
rect 56324 117215 56376 117224
rect 56324 117181 56333 117215
rect 56333 117181 56367 117215
rect 56367 117181 56376 117215
rect 56324 117172 56376 117181
rect 58624 117104 58676 117156
rect 66536 117104 66588 117156
rect 70860 117240 70912 117292
rect 67272 117147 67324 117156
rect 67272 117113 67281 117147
rect 67281 117113 67315 117147
rect 67315 117113 67324 117147
rect 67272 117104 67324 117113
rect 78588 117240 78640 117292
rect 77944 117172 77996 117224
rect 75000 117147 75052 117156
rect 75000 117113 75009 117147
rect 75009 117113 75043 117147
rect 75043 117113 75052 117147
rect 75000 117104 75052 117113
rect 41420 117036 41472 117088
rect 49056 117079 49108 117088
rect 49056 117045 49065 117079
rect 49065 117045 49099 117079
rect 49099 117045 49108 117079
rect 49056 117036 49108 117045
rect 64052 117079 64104 117088
rect 64052 117045 64061 117079
rect 64061 117045 64095 117079
rect 64095 117045 64104 117079
rect 64052 117036 64104 117045
rect 66720 117079 66772 117088
rect 66720 117045 66729 117079
rect 66729 117045 66763 117079
rect 66763 117045 66772 117079
rect 66720 117036 66772 117045
rect 71320 117079 71372 117088
rect 71320 117045 71329 117079
rect 71329 117045 71363 117079
rect 71363 117045 71372 117079
rect 71320 117036 71372 117045
rect 74540 117079 74592 117088
rect 74540 117045 74549 117079
rect 74549 117045 74583 117079
rect 74583 117045 74592 117079
rect 74540 117036 74592 117045
rect 4214 116934 4266 116986
rect 4278 116934 4330 116986
rect 4342 116934 4394 116986
rect 4406 116934 4458 116986
rect 4470 116934 4522 116986
rect 34934 116934 34986 116986
rect 34998 116934 35050 116986
rect 35062 116934 35114 116986
rect 35126 116934 35178 116986
rect 35190 116934 35242 116986
rect 65654 116934 65706 116986
rect 65718 116934 65770 116986
rect 65782 116934 65834 116986
rect 65846 116934 65898 116986
rect 65910 116934 65962 116986
rect 15568 116832 15620 116884
rect 40776 116832 40828 116884
rect 41420 116832 41472 116884
rect 66720 116832 66772 116884
rect 77208 116832 77260 116884
rect 10692 116764 10744 116816
rect 34704 116764 34756 116816
rect 40040 116696 40092 116748
rect 74540 116696 74592 116748
rect 1860 116671 1912 116680
rect 1860 116637 1869 116671
rect 1869 116637 1903 116671
rect 1903 116637 1912 116671
rect 1860 116628 1912 116637
rect 77852 116671 77904 116680
rect 77852 116637 77861 116671
rect 77861 116637 77895 116671
rect 77895 116637 77904 116671
rect 77852 116628 77904 116637
rect 2228 116603 2280 116612
rect 2228 116569 2237 116603
rect 2237 116569 2271 116603
rect 2271 116569 2280 116603
rect 2228 116560 2280 116569
rect 19574 116390 19626 116442
rect 19638 116390 19690 116442
rect 19702 116390 19754 116442
rect 19766 116390 19818 116442
rect 19830 116390 19882 116442
rect 50294 116390 50346 116442
rect 50358 116390 50410 116442
rect 50422 116390 50474 116442
rect 50486 116390 50538 116442
rect 50550 116390 50602 116442
rect 40776 116331 40828 116340
rect 40776 116297 40785 116331
rect 40785 116297 40819 116331
rect 40819 116297 40828 116331
rect 40776 116288 40828 116297
rect 37464 116152 37516 116204
rect 49056 116152 49108 116204
rect 77852 115948 77904 116000
rect 4214 115846 4266 115898
rect 4278 115846 4330 115898
rect 4342 115846 4394 115898
rect 4406 115846 4458 115898
rect 4470 115846 4522 115898
rect 34934 115846 34986 115898
rect 34998 115846 35050 115898
rect 35062 115846 35114 115898
rect 35126 115846 35178 115898
rect 35190 115846 35242 115898
rect 65654 115846 65706 115898
rect 65718 115846 65770 115898
rect 65782 115846 65834 115898
rect 65846 115846 65898 115898
rect 65910 115846 65962 115898
rect 19574 115302 19626 115354
rect 19638 115302 19690 115354
rect 19702 115302 19754 115354
rect 19766 115302 19818 115354
rect 19830 115302 19882 115354
rect 50294 115302 50346 115354
rect 50358 115302 50410 115354
rect 50422 115302 50474 115354
rect 50486 115302 50538 115354
rect 50550 115302 50602 115354
rect 4214 114758 4266 114810
rect 4278 114758 4330 114810
rect 4342 114758 4394 114810
rect 4406 114758 4458 114810
rect 4470 114758 4522 114810
rect 34934 114758 34986 114810
rect 34998 114758 35050 114810
rect 35062 114758 35114 114810
rect 35126 114758 35178 114810
rect 35190 114758 35242 114810
rect 65654 114758 65706 114810
rect 65718 114758 65770 114810
rect 65782 114758 65834 114810
rect 65846 114758 65898 114810
rect 65910 114758 65962 114810
rect 77392 114452 77444 114504
rect 78036 114359 78088 114368
rect 78036 114325 78045 114359
rect 78045 114325 78079 114359
rect 78079 114325 78088 114359
rect 78036 114316 78088 114325
rect 19574 114214 19626 114266
rect 19638 114214 19690 114266
rect 19702 114214 19754 114266
rect 19766 114214 19818 114266
rect 19830 114214 19882 114266
rect 50294 114214 50346 114266
rect 50358 114214 50410 114266
rect 50422 114214 50474 114266
rect 50486 114214 50538 114266
rect 50550 114214 50602 114266
rect 28264 114112 28316 114164
rect 20628 113976 20680 114028
rect 4214 113670 4266 113722
rect 4278 113670 4330 113722
rect 4342 113670 4394 113722
rect 4406 113670 4458 113722
rect 4470 113670 4522 113722
rect 34934 113670 34986 113722
rect 34998 113670 35050 113722
rect 35062 113670 35114 113722
rect 35126 113670 35178 113722
rect 35190 113670 35242 113722
rect 65654 113670 65706 113722
rect 65718 113670 65770 113722
rect 65782 113670 65834 113722
rect 65846 113670 65898 113722
rect 65910 113670 65962 113722
rect 1400 113407 1452 113416
rect 1400 113373 1409 113407
rect 1409 113373 1443 113407
rect 1443 113373 1452 113407
rect 1400 113364 1452 113373
rect 1584 113271 1636 113280
rect 1584 113237 1593 113271
rect 1593 113237 1627 113271
rect 1627 113237 1636 113271
rect 1584 113228 1636 113237
rect 19574 113126 19626 113178
rect 19638 113126 19690 113178
rect 19702 113126 19754 113178
rect 19766 113126 19818 113178
rect 19830 113126 19882 113178
rect 50294 113126 50346 113178
rect 50358 113126 50410 113178
rect 50422 113126 50474 113178
rect 50486 113126 50538 113178
rect 50550 113126 50602 113178
rect 4214 112582 4266 112634
rect 4278 112582 4330 112634
rect 4342 112582 4394 112634
rect 4406 112582 4458 112634
rect 4470 112582 4522 112634
rect 34934 112582 34986 112634
rect 34998 112582 35050 112634
rect 35062 112582 35114 112634
rect 35126 112582 35178 112634
rect 35190 112582 35242 112634
rect 65654 112582 65706 112634
rect 65718 112582 65770 112634
rect 65782 112582 65834 112634
rect 65846 112582 65898 112634
rect 65910 112582 65962 112634
rect 19574 112038 19626 112090
rect 19638 112038 19690 112090
rect 19702 112038 19754 112090
rect 19766 112038 19818 112090
rect 19830 112038 19882 112090
rect 50294 112038 50346 112090
rect 50358 112038 50410 112090
rect 50422 112038 50474 112090
rect 50486 112038 50538 112090
rect 50550 112038 50602 112090
rect 66536 111911 66588 111920
rect 66536 111877 66545 111911
rect 66545 111877 66579 111911
rect 66579 111877 66588 111911
rect 66536 111868 66588 111877
rect 76012 111800 76064 111852
rect 4214 111494 4266 111546
rect 4278 111494 4330 111546
rect 4342 111494 4394 111546
rect 4406 111494 4458 111546
rect 4470 111494 4522 111546
rect 34934 111494 34986 111546
rect 34998 111494 35050 111546
rect 35062 111494 35114 111546
rect 35126 111494 35178 111546
rect 35190 111494 35242 111546
rect 65654 111494 65706 111546
rect 65718 111494 65770 111546
rect 65782 111494 65834 111546
rect 65846 111494 65898 111546
rect 65910 111494 65962 111546
rect 19574 110950 19626 111002
rect 19638 110950 19690 111002
rect 19702 110950 19754 111002
rect 19766 110950 19818 111002
rect 19830 110950 19882 111002
rect 50294 110950 50346 111002
rect 50358 110950 50410 111002
rect 50422 110950 50474 111002
rect 50486 110950 50538 111002
rect 50550 110950 50602 111002
rect 77760 110712 77812 110764
rect 77852 110551 77904 110560
rect 77852 110517 77861 110551
rect 77861 110517 77895 110551
rect 77895 110517 77904 110551
rect 77852 110508 77904 110517
rect 4214 110406 4266 110458
rect 4278 110406 4330 110458
rect 4342 110406 4394 110458
rect 4406 110406 4458 110458
rect 4470 110406 4522 110458
rect 34934 110406 34986 110458
rect 34998 110406 35050 110458
rect 35062 110406 35114 110458
rect 35126 110406 35178 110458
rect 35190 110406 35242 110458
rect 65654 110406 65706 110458
rect 65718 110406 65770 110458
rect 65782 110406 65834 110458
rect 65846 110406 65898 110458
rect 65910 110406 65962 110458
rect 19574 109862 19626 109914
rect 19638 109862 19690 109914
rect 19702 109862 19754 109914
rect 19766 109862 19818 109914
rect 19830 109862 19882 109914
rect 50294 109862 50346 109914
rect 50358 109862 50410 109914
rect 50422 109862 50474 109914
rect 50486 109862 50538 109914
rect 50550 109862 50602 109914
rect 1860 109667 1912 109676
rect 1860 109633 1869 109667
rect 1869 109633 1903 109667
rect 1903 109633 1912 109667
rect 1860 109624 1912 109633
rect 20628 109420 20680 109472
rect 4214 109318 4266 109370
rect 4278 109318 4330 109370
rect 4342 109318 4394 109370
rect 4406 109318 4458 109370
rect 4470 109318 4522 109370
rect 34934 109318 34986 109370
rect 34998 109318 35050 109370
rect 35062 109318 35114 109370
rect 35126 109318 35178 109370
rect 35190 109318 35242 109370
rect 65654 109318 65706 109370
rect 65718 109318 65770 109370
rect 65782 109318 65834 109370
rect 65846 109318 65898 109370
rect 65910 109318 65962 109370
rect 40040 109259 40092 109268
rect 40040 109225 40049 109259
rect 40049 109225 40083 109259
rect 40083 109225 40092 109259
rect 40040 109216 40092 109225
rect 39856 109055 39908 109064
rect 39856 109021 39865 109055
rect 39865 109021 39899 109055
rect 39899 109021 39908 109055
rect 39856 109012 39908 109021
rect 19574 108774 19626 108826
rect 19638 108774 19690 108826
rect 19702 108774 19754 108826
rect 19766 108774 19818 108826
rect 19830 108774 19882 108826
rect 50294 108774 50346 108826
rect 50358 108774 50410 108826
rect 50422 108774 50474 108826
rect 50486 108774 50538 108826
rect 50550 108774 50602 108826
rect 4214 108230 4266 108282
rect 4278 108230 4330 108282
rect 4342 108230 4394 108282
rect 4406 108230 4458 108282
rect 4470 108230 4522 108282
rect 34934 108230 34986 108282
rect 34998 108230 35050 108282
rect 35062 108230 35114 108282
rect 35126 108230 35178 108282
rect 35190 108230 35242 108282
rect 65654 108230 65706 108282
rect 65718 108230 65770 108282
rect 65782 108230 65834 108282
rect 65846 108230 65898 108282
rect 65910 108230 65962 108282
rect 19574 107686 19626 107738
rect 19638 107686 19690 107738
rect 19702 107686 19754 107738
rect 19766 107686 19818 107738
rect 19830 107686 19882 107738
rect 50294 107686 50346 107738
rect 50358 107686 50410 107738
rect 50422 107686 50474 107738
rect 50486 107686 50538 107738
rect 50550 107686 50602 107738
rect 4214 107142 4266 107194
rect 4278 107142 4330 107194
rect 4342 107142 4394 107194
rect 4406 107142 4458 107194
rect 4470 107142 4522 107194
rect 34934 107142 34986 107194
rect 34998 107142 35050 107194
rect 35062 107142 35114 107194
rect 35126 107142 35178 107194
rect 35190 107142 35242 107194
rect 65654 107142 65706 107194
rect 65718 107142 65770 107194
rect 65782 107142 65834 107194
rect 65846 107142 65898 107194
rect 65910 107142 65962 107194
rect 19574 106598 19626 106650
rect 19638 106598 19690 106650
rect 19702 106598 19754 106650
rect 19766 106598 19818 106650
rect 19830 106598 19882 106650
rect 50294 106598 50346 106650
rect 50358 106598 50410 106650
rect 50422 106598 50474 106650
rect 50486 106598 50538 106650
rect 50550 106598 50602 106650
rect 76012 106360 76064 106412
rect 77852 106199 77904 106208
rect 77852 106165 77861 106199
rect 77861 106165 77895 106199
rect 77895 106165 77904 106199
rect 77852 106156 77904 106165
rect 4214 106054 4266 106106
rect 4278 106054 4330 106106
rect 4342 106054 4394 106106
rect 4406 106054 4458 106106
rect 4470 106054 4522 106106
rect 34934 106054 34986 106106
rect 34998 106054 35050 106106
rect 35062 106054 35114 106106
rect 35126 106054 35178 106106
rect 35190 106054 35242 106106
rect 65654 106054 65706 106106
rect 65718 106054 65770 106106
rect 65782 106054 65834 106106
rect 65846 106054 65898 106106
rect 65910 106054 65962 106106
rect 1400 105791 1452 105800
rect 1400 105757 1409 105791
rect 1409 105757 1443 105791
rect 1443 105757 1452 105791
rect 1400 105748 1452 105757
rect 1860 105680 1912 105732
rect 19574 105510 19626 105562
rect 19638 105510 19690 105562
rect 19702 105510 19754 105562
rect 19766 105510 19818 105562
rect 19830 105510 19882 105562
rect 50294 105510 50346 105562
rect 50358 105510 50410 105562
rect 50422 105510 50474 105562
rect 50486 105510 50538 105562
rect 50550 105510 50602 105562
rect 4214 104966 4266 105018
rect 4278 104966 4330 105018
rect 4342 104966 4394 105018
rect 4406 104966 4458 105018
rect 4470 104966 4522 105018
rect 34934 104966 34986 105018
rect 34998 104966 35050 105018
rect 35062 104966 35114 105018
rect 35126 104966 35178 105018
rect 35190 104966 35242 105018
rect 65654 104966 65706 105018
rect 65718 104966 65770 105018
rect 65782 104966 65834 105018
rect 65846 104966 65898 105018
rect 65910 104966 65962 105018
rect 19574 104422 19626 104474
rect 19638 104422 19690 104474
rect 19702 104422 19754 104474
rect 19766 104422 19818 104474
rect 19830 104422 19882 104474
rect 50294 104422 50346 104474
rect 50358 104422 50410 104474
rect 50422 104422 50474 104474
rect 50486 104422 50538 104474
rect 50550 104422 50602 104474
rect 4214 103878 4266 103930
rect 4278 103878 4330 103930
rect 4342 103878 4394 103930
rect 4406 103878 4458 103930
rect 4470 103878 4522 103930
rect 34934 103878 34986 103930
rect 34998 103878 35050 103930
rect 35062 103878 35114 103930
rect 35126 103878 35178 103930
rect 35190 103878 35242 103930
rect 65654 103878 65706 103930
rect 65718 103878 65770 103930
rect 65782 103878 65834 103930
rect 65846 103878 65898 103930
rect 65910 103878 65962 103930
rect 77944 103708 77996 103760
rect 78036 103615 78088 103624
rect 78036 103581 78045 103615
rect 78045 103581 78079 103615
rect 78079 103581 78088 103615
rect 78036 103572 78088 103581
rect 19574 103334 19626 103386
rect 19638 103334 19690 103386
rect 19702 103334 19754 103386
rect 19766 103334 19818 103386
rect 19830 103334 19882 103386
rect 50294 103334 50346 103386
rect 50358 103334 50410 103386
rect 50422 103334 50474 103386
rect 50486 103334 50538 103386
rect 50550 103334 50602 103386
rect 77300 103096 77352 103148
rect 77300 102935 77352 102944
rect 77300 102901 77309 102935
rect 77309 102901 77343 102935
rect 77343 102901 77352 102935
rect 77300 102892 77352 102901
rect 77852 102935 77904 102944
rect 77852 102901 77861 102935
rect 77861 102901 77895 102935
rect 77895 102901 77904 102935
rect 77852 102892 77904 102901
rect 4214 102790 4266 102842
rect 4278 102790 4330 102842
rect 4342 102790 4394 102842
rect 4406 102790 4458 102842
rect 4470 102790 4522 102842
rect 34934 102790 34986 102842
rect 34998 102790 35050 102842
rect 35062 102790 35114 102842
rect 35126 102790 35178 102842
rect 35190 102790 35242 102842
rect 65654 102790 65706 102842
rect 65718 102790 65770 102842
rect 65782 102790 65834 102842
rect 65846 102790 65898 102842
rect 65910 102790 65962 102842
rect 19574 102246 19626 102298
rect 19638 102246 19690 102298
rect 19702 102246 19754 102298
rect 19766 102246 19818 102298
rect 19830 102246 19882 102298
rect 50294 102246 50346 102298
rect 50358 102246 50410 102298
rect 50422 102246 50474 102298
rect 50486 102246 50538 102298
rect 50550 102246 50602 102298
rect 4214 101702 4266 101754
rect 4278 101702 4330 101754
rect 4342 101702 4394 101754
rect 4406 101702 4458 101754
rect 4470 101702 4522 101754
rect 34934 101702 34986 101754
rect 34998 101702 35050 101754
rect 35062 101702 35114 101754
rect 35126 101702 35178 101754
rect 35190 101702 35242 101754
rect 65654 101702 65706 101754
rect 65718 101702 65770 101754
rect 65782 101702 65834 101754
rect 65846 101702 65898 101754
rect 65910 101702 65962 101754
rect 1400 101439 1452 101448
rect 1400 101405 1409 101439
rect 1409 101405 1443 101439
rect 1443 101405 1452 101439
rect 1400 101396 1452 101405
rect 39856 101260 39908 101312
rect 19574 101158 19626 101210
rect 19638 101158 19690 101210
rect 19702 101158 19754 101210
rect 19766 101158 19818 101210
rect 19830 101158 19882 101210
rect 50294 101158 50346 101210
rect 50358 101158 50410 101210
rect 50422 101158 50474 101210
rect 50486 101158 50538 101210
rect 50550 101158 50602 101210
rect 4214 100614 4266 100666
rect 4278 100614 4330 100666
rect 4342 100614 4394 100666
rect 4406 100614 4458 100666
rect 4470 100614 4522 100666
rect 34934 100614 34986 100666
rect 34998 100614 35050 100666
rect 35062 100614 35114 100666
rect 35126 100614 35178 100666
rect 35190 100614 35242 100666
rect 65654 100614 65706 100666
rect 65718 100614 65770 100666
rect 65782 100614 65834 100666
rect 65846 100614 65898 100666
rect 65910 100614 65962 100666
rect 58624 100555 58676 100564
rect 58624 100521 58633 100555
rect 58633 100521 58667 100555
rect 58667 100521 58676 100555
rect 58624 100512 58676 100521
rect 58532 100283 58584 100292
rect 58532 100249 58541 100283
rect 58541 100249 58575 100283
rect 58575 100249 58584 100283
rect 58532 100240 58584 100249
rect 19574 100070 19626 100122
rect 19638 100070 19690 100122
rect 19702 100070 19754 100122
rect 19766 100070 19818 100122
rect 19830 100070 19882 100122
rect 50294 100070 50346 100122
rect 50358 100070 50410 100122
rect 50422 100070 50474 100122
rect 50486 100070 50538 100122
rect 50550 100070 50602 100122
rect 4214 99526 4266 99578
rect 4278 99526 4330 99578
rect 4342 99526 4394 99578
rect 4406 99526 4458 99578
rect 4470 99526 4522 99578
rect 34934 99526 34986 99578
rect 34998 99526 35050 99578
rect 35062 99526 35114 99578
rect 35126 99526 35178 99578
rect 35190 99526 35242 99578
rect 65654 99526 65706 99578
rect 65718 99526 65770 99578
rect 65782 99526 65834 99578
rect 65846 99526 65898 99578
rect 65910 99526 65962 99578
rect 19574 98982 19626 99034
rect 19638 98982 19690 99034
rect 19702 98982 19754 99034
rect 19766 98982 19818 99034
rect 19830 98982 19882 99034
rect 50294 98982 50346 99034
rect 50358 98982 50410 99034
rect 50422 98982 50474 99034
rect 50486 98982 50538 99034
rect 50550 98982 50602 99034
rect 78128 98744 78180 98796
rect 77852 98651 77904 98660
rect 77852 98617 77861 98651
rect 77861 98617 77895 98651
rect 77895 98617 77904 98651
rect 77852 98608 77904 98617
rect 4214 98438 4266 98490
rect 4278 98438 4330 98490
rect 4342 98438 4394 98490
rect 4406 98438 4458 98490
rect 4470 98438 4522 98490
rect 34934 98438 34986 98490
rect 34998 98438 35050 98490
rect 35062 98438 35114 98490
rect 35126 98438 35178 98490
rect 35190 98438 35242 98490
rect 65654 98438 65706 98490
rect 65718 98438 65770 98490
rect 65782 98438 65834 98490
rect 65846 98438 65898 98490
rect 65910 98438 65962 98490
rect 19574 97894 19626 97946
rect 19638 97894 19690 97946
rect 19702 97894 19754 97946
rect 19766 97894 19818 97946
rect 19830 97894 19882 97946
rect 50294 97894 50346 97946
rect 50358 97894 50410 97946
rect 50422 97894 50474 97946
rect 50486 97894 50538 97946
rect 50550 97894 50602 97946
rect 1400 97699 1452 97708
rect 1400 97665 1409 97699
rect 1409 97665 1443 97699
rect 1443 97665 1452 97699
rect 1400 97656 1452 97665
rect 1676 97631 1728 97640
rect 1676 97597 1685 97631
rect 1685 97597 1719 97631
rect 1719 97597 1728 97631
rect 1676 97588 1728 97597
rect 4214 97350 4266 97402
rect 4278 97350 4330 97402
rect 4342 97350 4394 97402
rect 4406 97350 4458 97402
rect 4470 97350 4522 97402
rect 34934 97350 34986 97402
rect 34998 97350 35050 97402
rect 35062 97350 35114 97402
rect 35126 97350 35178 97402
rect 35190 97350 35242 97402
rect 65654 97350 65706 97402
rect 65718 97350 65770 97402
rect 65782 97350 65834 97402
rect 65846 97350 65898 97402
rect 65910 97350 65962 97402
rect 19574 96806 19626 96858
rect 19638 96806 19690 96858
rect 19702 96806 19754 96858
rect 19766 96806 19818 96858
rect 19830 96806 19882 96858
rect 50294 96806 50346 96858
rect 50358 96806 50410 96858
rect 50422 96806 50474 96858
rect 50486 96806 50538 96858
rect 50550 96806 50602 96858
rect 4214 96262 4266 96314
rect 4278 96262 4330 96314
rect 4342 96262 4394 96314
rect 4406 96262 4458 96314
rect 4470 96262 4522 96314
rect 34934 96262 34986 96314
rect 34998 96262 35050 96314
rect 35062 96262 35114 96314
rect 35126 96262 35178 96314
rect 35190 96262 35242 96314
rect 65654 96262 65706 96314
rect 65718 96262 65770 96314
rect 65782 96262 65834 96314
rect 65846 96262 65898 96314
rect 65910 96262 65962 96314
rect 40316 95931 40368 95940
rect 40316 95897 40325 95931
rect 40325 95897 40359 95931
rect 40359 95897 40368 95931
rect 40316 95888 40368 95897
rect 1492 95820 1544 95872
rect 19574 95718 19626 95770
rect 19638 95718 19690 95770
rect 19702 95718 19754 95770
rect 19766 95718 19818 95770
rect 19830 95718 19882 95770
rect 50294 95718 50346 95770
rect 50358 95718 50410 95770
rect 50422 95718 50474 95770
rect 50486 95718 50538 95770
rect 50550 95718 50602 95770
rect 4214 95174 4266 95226
rect 4278 95174 4330 95226
rect 4342 95174 4394 95226
rect 4406 95174 4458 95226
rect 4470 95174 4522 95226
rect 34934 95174 34986 95226
rect 34998 95174 35050 95226
rect 35062 95174 35114 95226
rect 35126 95174 35178 95226
rect 35190 95174 35242 95226
rect 65654 95174 65706 95226
rect 65718 95174 65770 95226
rect 65782 95174 65834 95226
rect 65846 95174 65898 95226
rect 65910 95174 65962 95226
rect 77944 94868 77996 94920
rect 78036 94775 78088 94784
rect 78036 94741 78045 94775
rect 78045 94741 78079 94775
rect 78079 94741 78088 94775
rect 78036 94732 78088 94741
rect 19574 94630 19626 94682
rect 19638 94630 19690 94682
rect 19702 94630 19754 94682
rect 19766 94630 19818 94682
rect 19830 94630 19882 94682
rect 50294 94630 50346 94682
rect 50358 94630 50410 94682
rect 50422 94630 50474 94682
rect 50486 94630 50538 94682
rect 50550 94630 50602 94682
rect 2964 94392 3016 94444
rect 1584 94231 1636 94240
rect 1584 94197 1593 94231
rect 1593 94197 1627 94231
rect 1627 94197 1636 94231
rect 1584 94188 1636 94197
rect 4214 94086 4266 94138
rect 4278 94086 4330 94138
rect 4342 94086 4394 94138
rect 4406 94086 4458 94138
rect 4470 94086 4522 94138
rect 34934 94086 34986 94138
rect 34998 94086 35050 94138
rect 35062 94086 35114 94138
rect 35126 94086 35178 94138
rect 35190 94086 35242 94138
rect 65654 94086 65706 94138
rect 65718 94086 65770 94138
rect 65782 94086 65834 94138
rect 65846 94086 65898 94138
rect 65910 94086 65962 94138
rect 19574 93542 19626 93594
rect 19638 93542 19690 93594
rect 19702 93542 19754 93594
rect 19766 93542 19818 93594
rect 19830 93542 19882 93594
rect 50294 93542 50346 93594
rect 50358 93542 50410 93594
rect 50422 93542 50474 93594
rect 50486 93542 50538 93594
rect 50550 93542 50602 93594
rect 4214 92998 4266 93050
rect 4278 92998 4330 93050
rect 4342 92998 4394 93050
rect 4406 92998 4458 93050
rect 4470 92998 4522 93050
rect 34934 92998 34986 93050
rect 34998 92998 35050 93050
rect 35062 92998 35114 93050
rect 35126 92998 35178 93050
rect 35190 92998 35242 93050
rect 65654 92998 65706 93050
rect 65718 92998 65770 93050
rect 65782 92998 65834 93050
rect 65846 92998 65898 93050
rect 65910 92998 65962 93050
rect 19574 92454 19626 92506
rect 19638 92454 19690 92506
rect 19702 92454 19754 92506
rect 19766 92454 19818 92506
rect 19830 92454 19882 92506
rect 50294 92454 50346 92506
rect 50358 92454 50410 92506
rect 50422 92454 50474 92506
rect 50486 92454 50538 92506
rect 50550 92454 50602 92506
rect 41420 92395 41472 92404
rect 41420 92361 41429 92395
rect 41429 92361 41463 92395
rect 41463 92361 41472 92395
rect 41420 92352 41472 92361
rect 41052 92216 41104 92268
rect 4214 91910 4266 91962
rect 4278 91910 4330 91962
rect 4342 91910 4394 91962
rect 4406 91910 4458 91962
rect 4470 91910 4522 91962
rect 34934 91910 34986 91962
rect 34998 91910 35050 91962
rect 35062 91910 35114 91962
rect 35126 91910 35178 91962
rect 35190 91910 35242 91962
rect 65654 91910 65706 91962
rect 65718 91910 65770 91962
rect 65782 91910 65834 91962
rect 65846 91910 65898 91962
rect 65910 91910 65962 91962
rect 19574 91366 19626 91418
rect 19638 91366 19690 91418
rect 19702 91366 19754 91418
rect 19766 91366 19818 91418
rect 19830 91366 19882 91418
rect 50294 91366 50346 91418
rect 50358 91366 50410 91418
rect 50422 91366 50474 91418
rect 50486 91366 50538 91418
rect 50550 91366 50602 91418
rect 4214 90822 4266 90874
rect 4278 90822 4330 90874
rect 4342 90822 4394 90874
rect 4406 90822 4458 90874
rect 4470 90822 4522 90874
rect 34934 90822 34986 90874
rect 34998 90822 35050 90874
rect 35062 90822 35114 90874
rect 35126 90822 35178 90874
rect 35190 90822 35242 90874
rect 65654 90822 65706 90874
rect 65718 90822 65770 90874
rect 65782 90822 65834 90874
rect 65846 90822 65898 90874
rect 65910 90822 65962 90874
rect 77944 90491 77996 90500
rect 77944 90457 77953 90491
rect 77953 90457 77987 90491
rect 77987 90457 77996 90491
rect 77944 90448 77996 90457
rect 58532 90380 58584 90432
rect 19574 90278 19626 90330
rect 19638 90278 19690 90330
rect 19702 90278 19754 90330
rect 19766 90278 19818 90330
rect 19830 90278 19882 90330
rect 50294 90278 50346 90330
rect 50358 90278 50410 90330
rect 50422 90278 50474 90330
rect 50486 90278 50538 90330
rect 50550 90278 50602 90330
rect 1492 90083 1544 90092
rect 1492 90049 1501 90083
rect 1501 90049 1535 90083
rect 1535 90049 1544 90083
rect 1492 90040 1544 90049
rect 41052 89972 41104 90024
rect 4214 89734 4266 89786
rect 4278 89734 4330 89786
rect 4342 89734 4394 89786
rect 4406 89734 4458 89786
rect 4470 89734 4522 89786
rect 34934 89734 34986 89786
rect 34998 89734 35050 89786
rect 35062 89734 35114 89786
rect 35126 89734 35178 89786
rect 35190 89734 35242 89786
rect 65654 89734 65706 89786
rect 65718 89734 65770 89786
rect 65782 89734 65834 89786
rect 65846 89734 65898 89786
rect 65910 89734 65962 89786
rect 19574 89190 19626 89242
rect 19638 89190 19690 89242
rect 19702 89190 19754 89242
rect 19766 89190 19818 89242
rect 19830 89190 19882 89242
rect 50294 89190 50346 89242
rect 50358 89190 50410 89242
rect 50422 89190 50474 89242
rect 50486 89190 50538 89242
rect 50550 89190 50602 89242
rect 39948 88995 40000 89004
rect 39948 88961 39957 88995
rect 39957 88961 39991 88995
rect 39991 88961 40000 88995
rect 39948 88952 40000 88961
rect 7840 88748 7892 88800
rect 4214 88646 4266 88698
rect 4278 88646 4330 88698
rect 4342 88646 4394 88698
rect 4406 88646 4458 88698
rect 4470 88646 4522 88698
rect 34934 88646 34986 88698
rect 34998 88646 35050 88698
rect 35062 88646 35114 88698
rect 35126 88646 35178 88698
rect 35190 88646 35242 88698
rect 65654 88646 65706 88698
rect 65718 88646 65770 88698
rect 65782 88646 65834 88698
rect 65846 88646 65898 88698
rect 65910 88646 65962 88698
rect 19574 88102 19626 88154
rect 19638 88102 19690 88154
rect 19702 88102 19754 88154
rect 19766 88102 19818 88154
rect 19830 88102 19882 88154
rect 50294 88102 50346 88154
rect 50358 88102 50410 88154
rect 50422 88102 50474 88154
rect 50486 88102 50538 88154
rect 50550 88102 50602 88154
rect 4214 87558 4266 87610
rect 4278 87558 4330 87610
rect 4342 87558 4394 87610
rect 4406 87558 4458 87610
rect 4470 87558 4522 87610
rect 34934 87558 34986 87610
rect 34998 87558 35050 87610
rect 35062 87558 35114 87610
rect 35126 87558 35178 87610
rect 35190 87558 35242 87610
rect 65654 87558 65706 87610
rect 65718 87558 65770 87610
rect 65782 87558 65834 87610
rect 65846 87558 65898 87610
rect 65910 87558 65962 87610
rect 77944 87184 77996 87236
rect 40316 87116 40368 87168
rect 19574 87014 19626 87066
rect 19638 87014 19690 87066
rect 19702 87014 19754 87066
rect 19766 87014 19818 87066
rect 19830 87014 19882 87066
rect 50294 87014 50346 87066
rect 50358 87014 50410 87066
rect 50422 87014 50474 87066
rect 50486 87014 50538 87066
rect 50550 87014 50602 87066
rect 4214 86470 4266 86522
rect 4278 86470 4330 86522
rect 4342 86470 4394 86522
rect 4406 86470 4458 86522
rect 4470 86470 4522 86522
rect 34934 86470 34986 86522
rect 34998 86470 35050 86522
rect 35062 86470 35114 86522
rect 35126 86470 35178 86522
rect 35190 86470 35242 86522
rect 65654 86470 65706 86522
rect 65718 86470 65770 86522
rect 65782 86470 65834 86522
rect 65846 86470 65898 86522
rect 65910 86470 65962 86522
rect 2044 86164 2096 86216
rect 1584 86071 1636 86080
rect 1584 86037 1593 86071
rect 1593 86037 1627 86071
rect 1627 86037 1636 86071
rect 1584 86028 1636 86037
rect 19574 85926 19626 85978
rect 19638 85926 19690 85978
rect 19702 85926 19754 85978
rect 19766 85926 19818 85978
rect 19830 85926 19882 85978
rect 50294 85926 50346 85978
rect 50358 85926 50410 85978
rect 50422 85926 50474 85978
rect 50486 85926 50538 85978
rect 50550 85926 50602 85978
rect 4214 85382 4266 85434
rect 4278 85382 4330 85434
rect 4342 85382 4394 85434
rect 4406 85382 4458 85434
rect 4470 85382 4522 85434
rect 34934 85382 34986 85434
rect 34998 85382 35050 85434
rect 35062 85382 35114 85434
rect 35126 85382 35178 85434
rect 35190 85382 35242 85434
rect 65654 85382 65706 85434
rect 65718 85382 65770 85434
rect 65782 85382 65834 85434
rect 65846 85382 65898 85434
rect 65910 85382 65962 85434
rect 19574 84838 19626 84890
rect 19638 84838 19690 84890
rect 19702 84838 19754 84890
rect 19766 84838 19818 84890
rect 19830 84838 19882 84890
rect 50294 84838 50346 84890
rect 50358 84838 50410 84890
rect 50422 84838 50474 84890
rect 50486 84838 50538 84890
rect 50550 84838 50602 84890
rect 4214 84294 4266 84346
rect 4278 84294 4330 84346
rect 4342 84294 4394 84346
rect 4406 84294 4458 84346
rect 4470 84294 4522 84346
rect 34934 84294 34986 84346
rect 34998 84294 35050 84346
rect 35062 84294 35114 84346
rect 35126 84294 35178 84346
rect 35190 84294 35242 84346
rect 65654 84294 65706 84346
rect 65718 84294 65770 84346
rect 65782 84294 65834 84346
rect 65846 84294 65898 84346
rect 65910 84294 65962 84346
rect 19574 83750 19626 83802
rect 19638 83750 19690 83802
rect 19702 83750 19754 83802
rect 19766 83750 19818 83802
rect 19830 83750 19882 83802
rect 50294 83750 50346 83802
rect 50358 83750 50410 83802
rect 50422 83750 50474 83802
rect 50486 83750 50538 83802
rect 50550 83750 50602 83802
rect 77668 83555 77720 83564
rect 77668 83521 77677 83555
rect 77677 83521 77711 83555
rect 77711 83521 77720 83555
rect 77668 83512 77720 83521
rect 77852 83351 77904 83360
rect 77852 83317 77861 83351
rect 77861 83317 77895 83351
rect 77895 83317 77904 83351
rect 77852 83308 77904 83317
rect 4214 83206 4266 83258
rect 4278 83206 4330 83258
rect 4342 83206 4394 83258
rect 4406 83206 4458 83258
rect 4470 83206 4522 83258
rect 34934 83206 34986 83258
rect 34998 83206 35050 83258
rect 35062 83206 35114 83258
rect 35126 83206 35178 83258
rect 35190 83206 35242 83258
rect 65654 83206 65706 83258
rect 65718 83206 65770 83258
rect 65782 83206 65834 83258
rect 65846 83206 65898 83258
rect 65910 83206 65962 83258
rect 19574 82662 19626 82714
rect 19638 82662 19690 82714
rect 19702 82662 19754 82714
rect 19766 82662 19818 82714
rect 19830 82662 19882 82714
rect 50294 82662 50346 82714
rect 50358 82662 50410 82714
rect 50422 82662 50474 82714
rect 50486 82662 50538 82714
rect 50550 82662 50602 82714
rect 4214 82118 4266 82170
rect 4278 82118 4330 82170
rect 4342 82118 4394 82170
rect 4406 82118 4458 82170
rect 4470 82118 4522 82170
rect 34934 82118 34986 82170
rect 34998 82118 35050 82170
rect 35062 82118 35114 82170
rect 35126 82118 35178 82170
rect 35190 82118 35242 82170
rect 65654 82118 65706 82170
rect 65718 82118 65770 82170
rect 65782 82118 65834 82170
rect 65846 82118 65898 82170
rect 65910 82118 65962 82170
rect 1400 81855 1452 81864
rect 1400 81821 1409 81855
rect 1409 81821 1443 81855
rect 1443 81821 1452 81855
rect 1400 81812 1452 81821
rect 2136 81744 2188 81796
rect 19574 81574 19626 81626
rect 19638 81574 19690 81626
rect 19702 81574 19754 81626
rect 19766 81574 19818 81626
rect 19830 81574 19882 81626
rect 50294 81574 50346 81626
rect 50358 81574 50410 81626
rect 50422 81574 50474 81626
rect 50486 81574 50538 81626
rect 50550 81574 50602 81626
rect 4214 81030 4266 81082
rect 4278 81030 4330 81082
rect 4342 81030 4394 81082
rect 4406 81030 4458 81082
rect 4470 81030 4522 81082
rect 34934 81030 34986 81082
rect 34998 81030 35050 81082
rect 35062 81030 35114 81082
rect 35126 81030 35178 81082
rect 35190 81030 35242 81082
rect 65654 81030 65706 81082
rect 65718 81030 65770 81082
rect 65782 81030 65834 81082
rect 65846 81030 65898 81082
rect 65910 81030 65962 81082
rect 19574 80486 19626 80538
rect 19638 80486 19690 80538
rect 19702 80486 19754 80538
rect 19766 80486 19818 80538
rect 19830 80486 19882 80538
rect 50294 80486 50346 80538
rect 50358 80486 50410 80538
rect 50422 80486 50474 80538
rect 50486 80486 50538 80538
rect 50550 80486 50602 80538
rect 4214 79942 4266 79994
rect 4278 79942 4330 79994
rect 4342 79942 4394 79994
rect 4406 79942 4458 79994
rect 4470 79942 4522 79994
rect 34934 79942 34986 79994
rect 34998 79942 35050 79994
rect 35062 79942 35114 79994
rect 35126 79942 35178 79994
rect 35190 79942 35242 79994
rect 65654 79942 65706 79994
rect 65718 79942 65770 79994
rect 65782 79942 65834 79994
rect 65846 79942 65898 79994
rect 65910 79942 65962 79994
rect 19574 79398 19626 79450
rect 19638 79398 19690 79450
rect 19702 79398 19754 79450
rect 19766 79398 19818 79450
rect 19830 79398 19882 79450
rect 50294 79398 50346 79450
rect 50358 79398 50410 79450
rect 50422 79398 50474 79450
rect 50486 79398 50538 79450
rect 50550 79398 50602 79450
rect 10692 79339 10744 79348
rect 10692 79305 10701 79339
rect 10701 79305 10735 79339
rect 10735 79305 10744 79339
rect 10692 79296 10744 79305
rect 2780 79160 2832 79212
rect 77576 79203 77628 79212
rect 77576 79169 77585 79203
rect 77585 79169 77619 79203
rect 77619 79169 77628 79203
rect 77576 79160 77628 79169
rect 39948 78956 40000 79008
rect 4214 78854 4266 78906
rect 4278 78854 4330 78906
rect 4342 78854 4394 78906
rect 4406 78854 4458 78906
rect 4470 78854 4522 78906
rect 34934 78854 34986 78906
rect 34998 78854 35050 78906
rect 35062 78854 35114 78906
rect 35126 78854 35178 78906
rect 35190 78854 35242 78906
rect 65654 78854 65706 78906
rect 65718 78854 65770 78906
rect 65782 78854 65834 78906
rect 65846 78854 65898 78906
rect 65910 78854 65962 78906
rect 2596 78548 2648 78600
rect 1584 78455 1636 78464
rect 1584 78421 1593 78455
rect 1593 78421 1627 78455
rect 1627 78421 1636 78455
rect 1584 78412 1636 78421
rect 19574 78310 19626 78362
rect 19638 78310 19690 78362
rect 19702 78310 19754 78362
rect 19766 78310 19818 78362
rect 19830 78310 19882 78362
rect 50294 78310 50346 78362
rect 50358 78310 50410 78362
rect 50422 78310 50474 78362
rect 50486 78310 50538 78362
rect 50550 78310 50602 78362
rect 2596 78251 2648 78260
rect 2596 78217 2605 78251
rect 2605 78217 2639 78251
rect 2639 78217 2648 78251
rect 2596 78208 2648 78217
rect 2780 78115 2832 78124
rect 2780 78081 2789 78115
rect 2789 78081 2823 78115
rect 2823 78081 2832 78115
rect 2780 78072 2832 78081
rect 3056 78072 3108 78124
rect 4214 77766 4266 77818
rect 4278 77766 4330 77818
rect 4342 77766 4394 77818
rect 4406 77766 4458 77818
rect 4470 77766 4522 77818
rect 34934 77766 34986 77818
rect 34998 77766 35050 77818
rect 35062 77766 35114 77818
rect 35126 77766 35178 77818
rect 35190 77766 35242 77818
rect 65654 77766 65706 77818
rect 65718 77766 65770 77818
rect 65782 77766 65834 77818
rect 65846 77766 65898 77818
rect 65910 77766 65962 77818
rect 19574 77222 19626 77274
rect 19638 77222 19690 77274
rect 19702 77222 19754 77274
rect 19766 77222 19818 77274
rect 19830 77222 19882 77274
rect 50294 77222 50346 77274
rect 50358 77222 50410 77274
rect 50422 77222 50474 77274
rect 50486 77222 50538 77274
rect 50550 77222 50602 77274
rect 4214 76678 4266 76730
rect 4278 76678 4330 76730
rect 4342 76678 4394 76730
rect 4406 76678 4458 76730
rect 4470 76678 4522 76730
rect 34934 76678 34986 76730
rect 34998 76678 35050 76730
rect 35062 76678 35114 76730
rect 35126 76678 35178 76730
rect 35190 76678 35242 76730
rect 65654 76678 65706 76730
rect 65718 76678 65770 76730
rect 65782 76678 65834 76730
rect 65846 76678 65898 76730
rect 65910 76678 65962 76730
rect 19574 76134 19626 76186
rect 19638 76134 19690 76186
rect 19702 76134 19754 76186
rect 19766 76134 19818 76186
rect 19830 76134 19882 76186
rect 50294 76134 50346 76186
rect 50358 76134 50410 76186
rect 50422 76134 50474 76186
rect 50486 76134 50538 76186
rect 50550 76134 50602 76186
rect 4214 75590 4266 75642
rect 4278 75590 4330 75642
rect 4342 75590 4394 75642
rect 4406 75590 4458 75642
rect 4470 75590 4522 75642
rect 34934 75590 34986 75642
rect 34998 75590 35050 75642
rect 35062 75590 35114 75642
rect 35126 75590 35178 75642
rect 35190 75590 35242 75642
rect 65654 75590 65706 75642
rect 65718 75590 65770 75642
rect 65782 75590 65834 75642
rect 65846 75590 65898 75642
rect 65910 75590 65962 75642
rect 77944 75284 77996 75336
rect 78036 75191 78088 75200
rect 78036 75157 78045 75191
rect 78045 75157 78079 75191
rect 78079 75157 78088 75191
rect 78036 75148 78088 75157
rect 19574 75046 19626 75098
rect 19638 75046 19690 75098
rect 19702 75046 19754 75098
rect 19766 75046 19818 75098
rect 19830 75046 19882 75098
rect 50294 75046 50346 75098
rect 50358 75046 50410 75098
rect 50422 75046 50474 75098
rect 50486 75046 50538 75098
rect 50550 75046 50602 75098
rect 4214 74502 4266 74554
rect 4278 74502 4330 74554
rect 4342 74502 4394 74554
rect 4406 74502 4458 74554
rect 4470 74502 4522 74554
rect 34934 74502 34986 74554
rect 34998 74502 35050 74554
rect 35062 74502 35114 74554
rect 35126 74502 35178 74554
rect 35190 74502 35242 74554
rect 65654 74502 65706 74554
rect 65718 74502 65770 74554
rect 65782 74502 65834 74554
rect 65846 74502 65898 74554
rect 65910 74502 65962 74554
rect 1676 74264 1728 74316
rect 1952 74264 2004 74316
rect 1492 74196 1544 74248
rect 1584 74103 1636 74112
rect 1584 74069 1593 74103
rect 1593 74069 1627 74103
rect 1627 74069 1636 74103
rect 1584 74060 1636 74069
rect 19574 73958 19626 74010
rect 19638 73958 19690 74010
rect 19702 73958 19754 74010
rect 19766 73958 19818 74010
rect 19830 73958 19882 74010
rect 50294 73958 50346 74010
rect 50358 73958 50410 74010
rect 50422 73958 50474 74010
rect 50486 73958 50538 74010
rect 50550 73958 50602 74010
rect 4214 73414 4266 73466
rect 4278 73414 4330 73466
rect 4342 73414 4394 73466
rect 4406 73414 4458 73466
rect 4470 73414 4522 73466
rect 34934 73414 34986 73466
rect 34998 73414 35050 73466
rect 35062 73414 35114 73466
rect 35126 73414 35178 73466
rect 35190 73414 35242 73466
rect 65654 73414 65706 73466
rect 65718 73414 65770 73466
rect 65782 73414 65834 73466
rect 65846 73414 65898 73466
rect 65910 73414 65962 73466
rect 19574 72870 19626 72922
rect 19638 72870 19690 72922
rect 19702 72870 19754 72922
rect 19766 72870 19818 72922
rect 19830 72870 19882 72922
rect 50294 72870 50346 72922
rect 50358 72870 50410 72922
rect 50422 72870 50474 72922
rect 50486 72870 50538 72922
rect 50550 72870 50602 72922
rect 4214 72326 4266 72378
rect 4278 72326 4330 72378
rect 4342 72326 4394 72378
rect 4406 72326 4458 72378
rect 4470 72326 4522 72378
rect 34934 72326 34986 72378
rect 34998 72326 35050 72378
rect 35062 72326 35114 72378
rect 35126 72326 35178 72378
rect 35190 72326 35242 72378
rect 65654 72326 65706 72378
rect 65718 72326 65770 72378
rect 65782 72326 65834 72378
rect 65846 72326 65898 72378
rect 65910 72326 65962 72378
rect 76748 72020 76800 72072
rect 45192 71952 45244 72004
rect 19574 71782 19626 71834
rect 19638 71782 19690 71834
rect 19702 71782 19754 71834
rect 19766 71782 19818 71834
rect 19830 71782 19882 71834
rect 50294 71782 50346 71834
rect 50358 71782 50410 71834
rect 50422 71782 50474 71834
rect 50486 71782 50538 71834
rect 50550 71782 50602 71834
rect 76564 71544 76616 71596
rect 77852 71451 77904 71460
rect 77852 71417 77861 71451
rect 77861 71417 77895 71451
rect 77895 71417 77904 71451
rect 77852 71408 77904 71417
rect 4214 71238 4266 71290
rect 4278 71238 4330 71290
rect 4342 71238 4394 71290
rect 4406 71238 4458 71290
rect 4470 71238 4522 71290
rect 34934 71238 34986 71290
rect 34998 71238 35050 71290
rect 35062 71238 35114 71290
rect 35126 71238 35178 71290
rect 35190 71238 35242 71290
rect 65654 71238 65706 71290
rect 65718 71238 65770 71290
rect 65782 71238 65834 71290
rect 65846 71238 65898 71290
rect 65910 71238 65962 71290
rect 76564 71179 76616 71188
rect 76564 71145 76573 71179
rect 76573 71145 76607 71179
rect 76607 71145 76616 71179
rect 76564 71136 76616 71145
rect 2044 71111 2096 71120
rect 2044 71077 2053 71111
rect 2053 71077 2087 71111
rect 2087 71077 2096 71111
rect 2044 71068 2096 71077
rect 76748 70975 76800 70984
rect 76748 70941 76757 70975
rect 76757 70941 76791 70975
rect 76791 70941 76800 70975
rect 76748 70932 76800 70941
rect 77668 70932 77720 70984
rect 1676 70864 1728 70916
rect 19574 70694 19626 70746
rect 19638 70694 19690 70746
rect 19702 70694 19754 70746
rect 19766 70694 19818 70746
rect 19830 70694 19882 70746
rect 50294 70694 50346 70746
rect 50358 70694 50410 70746
rect 50422 70694 50474 70746
rect 50486 70694 50538 70746
rect 50550 70694 50602 70746
rect 1400 70499 1452 70508
rect 1400 70465 1409 70499
rect 1409 70465 1443 70499
rect 1443 70465 1452 70499
rect 1400 70456 1452 70465
rect 1584 70295 1636 70304
rect 1584 70261 1593 70295
rect 1593 70261 1627 70295
rect 1627 70261 1636 70295
rect 1584 70252 1636 70261
rect 4214 70150 4266 70202
rect 4278 70150 4330 70202
rect 4342 70150 4394 70202
rect 4406 70150 4458 70202
rect 4470 70150 4522 70202
rect 34934 70150 34986 70202
rect 34998 70150 35050 70202
rect 35062 70150 35114 70202
rect 35126 70150 35178 70202
rect 35190 70150 35242 70202
rect 65654 70150 65706 70202
rect 65718 70150 65770 70202
rect 65782 70150 65834 70202
rect 65846 70150 65898 70202
rect 65910 70150 65962 70202
rect 1400 70048 1452 70100
rect 1676 69844 1728 69896
rect 77484 69708 77536 69760
rect 77944 69708 77996 69760
rect 19574 69606 19626 69658
rect 19638 69606 19690 69658
rect 19702 69606 19754 69658
rect 19766 69606 19818 69658
rect 19830 69606 19882 69658
rect 50294 69606 50346 69658
rect 50358 69606 50410 69658
rect 50422 69606 50474 69658
rect 50486 69606 50538 69658
rect 50550 69606 50602 69658
rect 4214 69062 4266 69114
rect 4278 69062 4330 69114
rect 4342 69062 4394 69114
rect 4406 69062 4458 69114
rect 4470 69062 4522 69114
rect 34934 69062 34986 69114
rect 34998 69062 35050 69114
rect 35062 69062 35114 69114
rect 35126 69062 35178 69114
rect 35190 69062 35242 69114
rect 65654 69062 65706 69114
rect 65718 69062 65770 69114
rect 65782 69062 65834 69114
rect 65846 69062 65898 69114
rect 65910 69062 65962 69114
rect 19574 68518 19626 68570
rect 19638 68518 19690 68570
rect 19702 68518 19754 68570
rect 19766 68518 19818 68570
rect 19830 68518 19882 68570
rect 50294 68518 50346 68570
rect 50358 68518 50410 68570
rect 50422 68518 50474 68570
rect 50486 68518 50538 68570
rect 50550 68518 50602 68570
rect 4214 67974 4266 68026
rect 4278 67974 4330 68026
rect 4342 67974 4394 68026
rect 4406 67974 4458 68026
rect 4470 67974 4522 68026
rect 34934 67974 34986 68026
rect 34998 67974 35050 68026
rect 35062 67974 35114 68026
rect 35126 67974 35178 68026
rect 35190 67974 35242 68026
rect 65654 67974 65706 68026
rect 65718 67974 65770 68026
rect 65782 67974 65834 68026
rect 65846 67974 65898 68026
rect 65910 67974 65962 68026
rect 77944 67600 77996 67652
rect 77852 67575 77904 67584
rect 77852 67541 77861 67575
rect 77861 67541 77895 67575
rect 77895 67541 77904 67575
rect 77852 67532 77904 67541
rect 19574 67430 19626 67482
rect 19638 67430 19690 67482
rect 19702 67430 19754 67482
rect 19766 67430 19818 67482
rect 19830 67430 19882 67482
rect 50294 67430 50346 67482
rect 50358 67430 50410 67482
rect 50422 67430 50474 67482
rect 50486 67430 50538 67482
rect 50550 67430 50602 67482
rect 4214 66886 4266 66938
rect 4278 66886 4330 66938
rect 4342 66886 4394 66938
rect 4406 66886 4458 66938
rect 4470 66886 4522 66938
rect 34934 66886 34986 66938
rect 34998 66886 35050 66938
rect 35062 66886 35114 66938
rect 35126 66886 35178 66938
rect 35190 66886 35242 66938
rect 65654 66886 65706 66938
rect 65718 66886 65770 66938
rect 65782 66886 65834 66938
rect 65846 66886 65898 66938
rect 65910 66886 65962 66938
rect 19574 66342 19626 66394
rect 19638 66342 19690 66394
rect 19702 66342 19754 66394
rect 19766 66342 19818 66394
rect 19830 66342 19882 66394
rect 50294 66342 50346 66394
rect 50358 66342 50410 66394
rect 50422 66342 50474 66394
rect 50486 66342 50538 66394
rect 50550 66342 50602 66394
rect 2320 66147 2372 66156
rect 1584 66011 1636 66020
rect 1584 65977 1593 66011
rect 1593 65977 1627 66011
rect 1627 65977 1636 66011
rect 1584 65968 1636 65977
rect 2320 66113 2329 66147
rect 2329 66113 2363 66147
rect 2363 66113 2372 66147
rect 2320 66104 2372 66113
rect 4214 65798 4266 65850
rect 4278 65798 4330 65850
rect 4342 65798 4394 65850
rect 4406 65798 4458 65850
rect 4470 65798 4522 65850
rect 34934 65798 34986 65850
rect 34998 65798 35050 65850
rect 35062 65798 35114 65850
rect 35126 65798 35178 65850
rect 35190 65798 35242 65850
rect 65654 65798 65706 65850
rect 65718 65798 65770 65850
rect 65782 65798 65834 65850
rect 65846 65798 65898 65850
rect 65910 65798 65962 65850
rect 40684 65560 40736 65612
rect 2320 65492 2372 65544
rect 39856 65535 39908 65544
rect 39856 65501 39865 65535
rect 39865 65501 39899 65535
rect 39899 65501 39908 65535
rect 39856 65492 39908 65501
rect 11888 65424 11940 65476
rect 1768 65356 1820 65408
rect 40040 65424 40092 65476
rect 19574 65254 19626 65306
rect 19638 65254 19690 65306
rect 19702 65254 19754 65306
rect 19766 65254 19818 65306
rect 19830 65254 19882 65306
rect 50294 65254 50346 65306
rect 50358 65254 50410 65306
rect 50422 65254 50474 65306
rect 50486 65254 50538 65306
rect 50550 65254 50602 65306
rect 40040 65195 40092 65204
rect 40040 65161 40049 65195
rect 40049 65161 40083 65195
rect 40083 65161 40092 65195
rect 40040 65152 40092 65161
rect 41052 65195 41104 65204
rect 41052 65161 41061 65195
rect 41061 65161 41095 65195
rect 41095 65161 41104 65195
rect 41052 65152 41104 65161
rect 40684 64991 40736 65000
rect 40684 64957 40693 64991
rect 40693 64957 40727 64991
rect 40727 64957 40736 64991
rect 40684 64948 40736 64957
rect 40868 64812 40920 64864
rect 41696 64812 41748 64864
rect 77852 64812 77904 64864
rect 4214 64710 4266 64762
rect 4278 64710 4330 64762
rect 4342 64710 4394 64762
rect 4406 64710 4458 64762
rect 4470 64710 4522 64762
rect 34934 64710 34986 64762
rect 34998 64710 35050 64762
rect 35062 64710 35114 64762
rect 35126 64710 35178 64762
rect 35190 64710 35242 64762
rect 65654 64710 65706 64762
rect 65718 64710 65770 64762
rect 65782 64710 65834 64762
rect 65846 64710 65898 64762
rect 65910 64710 65962 64762
rect 39488 64404 39540 64456
rect 41696 64540 41748 64592
rect 40500 64447 40552 64456
rect 40500 64413 40509 64447
rect 40509 64413 40543 64447
rect 40543 64413 40552 64447
rect 40500 64404 40552 64413
rect 41052 64472 41104 64524
rect 40868 64447 40920 64456
rect 40868 64413 40877 64447
rect 40877 64413 40911 64447
rect 40911 64413 40920 64447
rect 40868 64404 40920 64413
rect 19574 64166 19626 64218
rect 19638 64166 19690 64218
rect 19702 64166 19754 64218
rect 19766 64166 19818 64218
rect 19830 64166 19882 64218
rect 50294 64166 50346 64218
rect 50358 64166 50410 64218
rect 50422 64166 50474 64218
rect 50486 64166 50538 64218
rect 50550 64166 50602 64218
rect 39488 63971 39540 63980
rect 39488 63937 39497 63971
rect 39497 63937 39531 63971
rect 39531 63937 39540 63971
rect 39488 63928 39540 63937
rect 39488 63724 39540 63776
rect 4214 63622 4266 63674
rect 4278 63622 4330 63674
rect 4342 63622 4394 63674
rect 4406 63622 4458 63674
rect 4470 63622 4522 63674
rect 34934 63622 34986 63674
rect 34998 63622 35050 63674
rect 35062 63622 35114 63674
rect 35126 63622 35178 63674
rect 35190 63622 35242 63674
rect 65654 63622 65706 63674
rect 65718 63622 65770 63674
rect 65782 63622 65834 63674
rect 65846 63622 65898 63674
rect 65910 63622 65962 63674
rect 38292 63316 38344 63368
rect 78036 63223 78088 63232
rect 78036 63189 78045 63223
rect 78045 63189 78079 63223
rect 78079 63189 78088 63223
rect 78036 63180 78088 63189
rect 19574 63078 19626 63130
rect 19638 63078 19690 63130
rect 19702 63078 19754 63130
rect 19766 63078 19818 63130
rect 19830 63078 19882 63130
rect 50294 63078 50346 63130
rect 50358 63078 50410 63130
rect 50422 63078 50474 63130
rect 50486 63078 50538 63130
rect 50550 63078 50602 63130
rect 1400 62883 1452 62892
rect 1400 62849 1409 62883
rect 1409 62849 1443 62883
rect 1443 62849 1452 62883
rect 1400 62840 1452 62849
rect 1584 62679 1636 62688
rect 1584 62645 1593 62679
rect 1593 62645 1627 62679
rect 1627 62645 1636 62679
rect 1584 62636 1636 62645
rect 4214 62534 4266 62586
rect 4278 62534 4330 62586
rect 4342 62534 4394 62586
rect 4406 62534 4458 62586
rect 4470 62534 4522 62586
rect 34934 62534 34986 62586
rect 34998 62534 35050 62586
rect 35062 62534 35114 62586
rect 35126 62534 35178 62586
rect 35190 62534 35242 62586
rect 65654 62534 65706 62586
rect 65718 62534 65770 62586
rect 65782 62534 65834 62586
rect 65846 62534 65898 62586
rect 65910 62534 65962 62586
rect 19574 61990 19626 62042
rect 19638 61990 19690 62042
rect 19702 61990 19754 62042
rect 19766 61990 19818 62042
rect 19830 61990 19882 62042
rect 50294 61990 50346 62042
rect 50358 61990 50410 62042
rect 50422 61990 50474 62042
rect 50486 61990 50538 62042
rect 50550 61990 50602 62042
rect 4214 61446 4266 61498
rect 4278 61446 4330 61498
rect 4342 61446 4394 61498
rect 4406 61446 4458 61498
rect 4470 61446 4522 61498
rect 34934 61446 34986 61498
rect 34998 61446 35050 61498
rect 35062 61446 35114 61498
rect 35126 61446 35178 61498
rect 35190 61446 35242 61498
rect 65654 61446 65706 61498
rect 65718 61446 65770 61498
rect 65782 61446 65834 61498
rect 65846 61446 65898 61498
rect 65910 61446 65962 61498
rect 39764 61140 39816 61192
rect 19432 61072 19484 61124
rect 19574 60902 19626 60954
rect 19638 60902 19690 60954
rect 19702 60902 19754 60954
rect 19766 60902 19818 60954
rect 19830 60902 19882 60954
rect 50294 60902 50346 60954
rect 50358 60902 50410 60954
rect 50422 60902 50474 60954
rect 50486 60902 50538 60954
rect 50550 60902 50602 60954
rect 39948 60775 40000 60784
rect 39948 60741 39957 60775
rect 39957 60741 39991 60775
rect 39991 60741 40000 60775
rect 39948 60732 40000 60741
rect 40776 60732 40828 60784
rect 38844 60664 38896 60716
rect 77300 60596 77352 60648
rect 1492 60528 1544 60580
rect 77576 60460 77628 60512
rect 4214 60358 4266 60410
rect 4278 60358 4330 60410
rect 4342 60358 4394 60410
rect 4406 60358 4458 60410
rect 4470 60358 4522 60410
rect 34934 60358 34986 60410
rect 34998 60358 35050 60410
rect 35062 60358 35114 60410
rect 35126 60358 35178 60410
rect 35190 60358 35242 60410
rect 65654 60358 65706 60410
rect 65718 60358 65770 60410
rect 65782 60358 65834 60410
rect 65846 60358 65898 60410
rect 65910 60358 65962 60410
rect 2136 60256 2188 60308
rect 35808 60299 35860 60308
rect 1860 60120 1912 60172
rect 35808 60265 35817 60299
rect 35817 60265 35851 60299
rect 35851 60265 35860 60299
rect 35808 60256 35860 60265
rect 36360 60299 36412 60308
rect 36360 60265 36369 60299
rect 36369 60265 36403 60299
rect 36403 60265 36412 60299
rect 36360 60256 36412 60265
rect 38292 60299 38344 60308
rect 38292 60265 38301 60299
rect 38301 60265 38335 60299
rect 38335 60265 38344 60299
rect 38292 60256 38344 60265
rect 77760 60256 77812 60308
rect 2228 60052 2280 60104
rect 22652 60120 22704 60172
rect 41052 60095 41104 60104
rect 19984 59984 20036 60036
rect 35808 59984 35860 60036
rect 36268 60027 36320 60036
rect 36268 59993 36277 60027
rect 36277 59993 36311 60027
rect 36311 59993 36320 60027
rect 36268 59984 36320 59993
rect 41052 60061 41061 60095
rect 41061 60061 41095 60095
rect 41095 60061 41104 60095
rect 41052 60052 41104 60061
rect 56324 60052 56376 60104
rect 38936 60027 38988 60036
rect 38936 59993 38945 60027
rect 38945 59993 38979 60027
rect 38979 59993 38988 60027
rect 38936 59984 38988 59993
rect 40592 59984 40644 60036
rect 77760 60027 77812 60036
rect 1492 59916 1544 59968
rect 35348 59916 35400 59968
rect 37740 59959 37792 59968
rect 37740 59925 37749 59959
rect 37749 59925 37783 59959
rect 37783 59925 37792 59959
rect 37740 59916 37792 59925
rect 63040 59959 63092 59968
rect 63040 59925 63049 59959
rect 63049 59925 63083 59959
rect 63083 59925 63092 59959
rect 63040 59916 63092 59925
rect 77760 59993 77769 60027
rect 77769 59993 77803 60027
rect 77803 59993 77812 60027
rect 77760 59984 77812 59993
rect 77484 59916 77536 59968
rect 19574 59814 19626 59866
rect 19638 59814 19690 59866
rect 19702 59814 19754 59866
rect 19766 59814 19818 59866
rect 19830 59814 19882 59866
rect 50294 59814 50346 59866
rect 50358 59814 50410 59866
rect 50422 59814 50474 59866
rect 50486 59814 50538 59866
rect 50550 59814 50602 59866
rect 4620 59712 4672 59764
rect 33140 59712 33192 59764
rect 36268 59712 36320 59764
rect 77760 59755 77812 59764
rect 77760 59721 77769 59755
rect 77769 59721 77803 59755
rect 77803 59721 77812 59755
rect 77760 59712 77812 59721
rect 37740 59644 37792 59696
rect 1952 59576 2004 59628
rect 39580 59576 39632 59628
rect 41144 59576 41196 59628
rect 71320 59576 71372 59628
rect 77944 59619 77996 59628
rect 77944 59585 77953 59619
rect 77953 59585 77987 59619
rect 77987 59585 77996 59619
rect 77944 59576 77996 59585
rect 39120 59551 39172 59560
rect 39120 59517 39129 59551
rect 39129 59517 39163 59551
rect 39163 59517 39172 59551
rect 39120 59508 39172 59517
rect 77392 59508 77444 59560
rect 1400 59372 1452 59424
rect 77392 59372 77444 59424
rect 4214 59270 4266 59322
rect 4278 59270 4330 59322
rect 4342 59270 4394 59322
rect 4406 59270 4458 59322
rect 4470 59270 4522 59322
rect 34934 59270 34986 59322
rect 34998 59270 35050 59322
rect 35062 59270 35114 59322
rect 35126 59270 35178 59322
rect 35190 59270 35242 59322
rect 65654 59270 65706 59322
rect 65718 59270 65770 59322
rect 65782 59270 65834 59322
rect 65846 59270 65898 59322
rect 65910 59270 65962 59322
rect 2964 59211 3016 59220
rect 2964 59177 2973 59211
rect 2973 59177 3007 59211
rect 3007 59177 3016 59211
rect 2964 59168 3016 59177
rect 1400 59007 1452 59016
rect 1400 58973 1409 59007
rect 1409 58973 1443 59007
rect 1443 58973 1452 59007
rect 1400 58964 1452 58973
rect 2964 58964 3016 59016
rect 39672 58964 39724 59016
rect 63868 58896 63920 58948
rect 1584 58871 1636 58880
rect 1584 58837 1593 58871
rect 1593 58837 1627 58871
rect 1627 58837 1636 58871
rect 1584 58828 1636 58837
rect 19574 58726 19626 58778
rect 19638 58726 19690 58778
rect 19702 58726 19754 58778
rect 19766 58726 19818 58778
rect 19830 58726 19882 58778
rect 50294 58726 50346 58778
rect 50358 58726 50410 58778
rect 50422 58726 50474 58778
rect 50486 58726 50538 58778
rect 50550 58726 50602 58778
rect 1400 58624 1452 58676
rect 1676 58488 1728 58540
rect 2964 58531 3016 58540
rect 2964 58497 2973 58531
rect 2973 58497 3007 58531
rect 3007 58497 3016 58531
rect 2964 58488 3016 58497
rect 1676 58284 1728 58336
rect 4214 58182 4266 58234
rect 4278 58182 4330 58234
rect 4342 58182 4394 58234
rect 4406 58182 4458 58234
rect 4470 58182 4522 58234
rect 34934 58182 34986 58234
rect 34998 58182 35050 58234
rect 35062 58182 35114 58234
rect 35126 58182 35178 58234
rect 35190 58182 35242 58234
rect 65654 58182 65706 58234
rect 65718 58182 65770 58234
rect 65782 58182 65834 58234
rect 65846 58182 65898 58234
rect 65910 58182 65962 58234
rect 19574 57638 19626 57690
rect 19638 57638 19690 57690
rect 19702 57638 19754 57690
rect 19766 57638 19818 57690
rect 19830 57638 19882 57690
rect 50294 57638 50346 57690
rect 50358 57638 50410 57690
rect 50422 57638 50474 57690
rect 50486 57638 50538 57690
rect 50550 57638 50602 57690
rect 4214 57094 4266 57146
rect 4278 57094 4330 57146
rect 4342 57094 4394 57146
rect 4406 57094 4458 57146
rect 4470 57094 4522 57146
rect 34934 57094 34986 57146
rect 34998 57094 35050 57146
rect 35062 57094 35114 57146
rect 35126 57094 35178 57146
rect 35190 57094 35242 57146
rect 65654 57094 65706 57146
rect 65718 57094 65770 57146
rect 65782 57094 65834 57146
rect 65846 57094 65898 57146
rect 65910 57094 65962 57146
rect 19574 56550 19626 56602
rect 19638 56550 19690 56602
rect 19702 56550 19754 56602
rect 19766 56550 19818 56602
rect 19830 56550 19882 56602
rect 50294 56550 50346 56602
rect 50358 56550 50410 56602
rect 50422 56550 50474 56602
rect 50486 56550 50538 56602
rect 50550 56550 50602 56602
rect 77760 56312 77812 56364
rect 77852 56151 77904 56160
rect 77852 56117 77861 56151
rect 77861 56117 77895 56151
rect 77895 56117 77904 56151
rect 77852 56108 77904 56117
rect 4214 56006 4266 56058
rect 4278 56006 4330 56058
rect 4342 56006 4394 56058
rect 4406 56006 4458 56058
rect 4470 56006 4522 56058
rect 34934 56006 34986 56058
rect 34998 56006 35050 56058
rect 35062 56006 35114 56058
rect 35126 56006 35178 56058
rect 35190 56006 35242 56058
rect 65654 56006 65706 56058
rect 65718 56006 65770 56058
rect 65782 56006 65834 56058
rect 65846 56006 65898 56058
rect 65910 56006 65962 56058
rect 19574 55462 19626 55514
rect 19638 55462 19690 55514
rect 19702 55462 19754 55514
rect 19766 55462 19818 55514
rect 19830 55462 19882 55514
rect 50294 55462 50346 55514
rect 50358 55462 50410 55514
rect 50422 55462 50474 55514
rect 50486 55462 50538 55514
rect 50550 55462 50602 55514
rect 4214 54918 4266 54970
rect 4278 54918 4330 54970
rect 4342 54918 4394 54970
rect 4406 54918 4458 54970
rect 4470 54918 4522 54970
rect 34934 54918 34986 54970
rect 34998 54918 35050 54970
rect 35062 54918 35114 54970
rect 35126 54918 35178 54970
rect 35190 54918 35242 54970
rect 65654 54918 65706 54970
rect 65718 54918 65770 54970
rect 65782 54918 65834 54970
rect 65846 54918 65898 54970
rect 65910 54918 65962 54970
rect 40500 54612 40552 54664
rect 1492 54519 1544 54528
rect 1492 54485 1501 54519
rect 1501 54485 1535 54519
rect 1535 54485 1544 54519
rect 1492 54476 1544 54485
rect 19574 54374 19626 54426
rect 19638 54374 19690 54426
rect 19702 54374 19754 54426
rect 19766 54374 19818 54426
rect 19830 54374 19882 54426
rect 50294 54374 50346 54426
rect 50358 54374 50410 54426
rect 50422 54374 50474 54426
rect 50486 54374 50538 54426
rect 50550 54374 50602 54426
rect 4214 53830 4266 53882
rect 4278 53830 4330 53882
rect 4342 53830 4394 53882
rect 4406 53830 4458 53882
rect 4470 53830 4522 53882
rect 34934 53830 34986 53882
rect 34998 53830 35050 53882
rect 35062 53830 35114 53882
rect 35126 53830 35178 53882
rect 35190 53830 35242 53882
rect 65654 53830 65706 53882
rect 65718 53830 65770 53882
rect 65782 53830 65834 53882
rect 65846 53830 65898 53882
rect 65910 53830 65962 53882
rect 19574 53286 19626 53338
rect 19638 53286 19690 53338
rect 19702 53286 19754 53338
rect 19766 53286 19818 53338
rect 19830 53286 19882 53338
rect 50294 53286 50346 53338
rect 50358 53286 50410 53338
rect 50422 53286 50474 53338
rect 50486 53286 50538 53338
rect 50550 53286 50602 53338
rect 4214 52742 4266 52794
rect 4278 52742 4330 52794
rect 4342 52742 4394 52794
rect 4406 52742 4458 52794
rect 4470 52742 4522 52794
rect 34934 52742 34986 52794
rect 34998 52742 35050 52794
rect 35062 52742 35114 52794
rect 35126 52742 35178 52794
rect 35190 52742 35242 52794
rect 65654 52742 65706 52794
rect 65718 52742 65770 52794
rect 65782 52742 65834 52794
rect 65846 52742 65898 52794
rect 65910 52742 65962 52794
rect 19574 52198 19626 52250
rect 19638 52198 19690 52250
rect 19702 52198 19754 52250
rect 19766 52198 19818 52250
rect 19830 52198 19882 52250
rect 50294 52198 50346 52250
rect 50358 52198 50410 52250
rect 50422 52198 50474 52250
rect 50486 52198 50538 52250
rect 50550 52198 50602 52250
rect 77392 51960 77444 52012
rect 77852 51799 77904 51808
rect 77852 51765 77861 51799
rect 77861 51765 77895 51799
rect 77895 51765 77904 51799
rect 77852 51756 77904 51765
rect 4214 51654 4266 51706
rect 4278 51654 4330 51706
rect 4342 51654 4394 51706
rect 4406 51654 4458 51706
rect 4470 51654 4522 51706
rect 34934 51654 34986 51706
rect 34998 51654 35050 51706
rect 35062 51654 35114 51706
rect 35126 51654 35178 51706
rect 35190 51654 35242 51706
rect 65654 51654 65706 51706
rect 65718 51654 65770 51706
rect 65782 51654 65834 51706
rect 65846 51654 65898 51706
rect 65910 51654 65962 51706
rect 19574 51110 19626 51162
rect 19638 51110 19690 51162
rect 19702 51110 19754 51162
rect 19766 51110 19818 51162
rect 19830 51110 19882 51162
rect 50294 51110 50346 51162
rect 50358 51110 50410 51162
rect 50422 51110 50474 51162
rect 50486 51110 50538 51162
rect 50550 51110 50602 51162
rect 39488 50872 39540 50924
rect 1492 50711 1544 50720
rect 1492 50677 1501 50711
rect 1501 50677 1535 50711
rect 1535 50677 1544 50711
rect 1492 50668 1544 50677
rect 4214 50566 4266 50618
rect 4278 50566 4330 50618
rect 4342 50566 4394 50618
rect 4406 50566 4458 50618
rect 4470 50566 4522 50618
rect 34934 50566 34986 50618
rect 34998 50566 35050 50618
rect 35062 50566 35114 50618
rect 35126 50566 35178 50618
rect 35190 50566 35242 50618
rect 65654 50566 65706 50618
rect 65718 50566 65770 50618
rect 65782 50566 65834 50618
rect 65846 50566 65898 50618
rect 65910 50566 65962 50618
rect 19574 50022 19626 50074
rect 19638 50022 19690 50074
rect 19702 50022 19754 50074
rect 19766 50022 19818 50074
rect 19830 50022 19882 50074
rect 50294 50022 50346 50074
rect 50358 50022 50410 50074
rect 50422 50022 50474 50074
rect 50486 50022 50538 50074
rect 50550 50022 50602 50074
rect 4214 49478 4266 49530
rect 4278 49478 4330 49530
rect 4342 49478 4394 49530
rect 4406 49478 4458 49530
rect 4470 49478 4522 49530
rect 34934 49478 34986 49530
rect 34998 49478 35050 49530
rect 35062 49478 35114 49530
rect 35126 49478 35178 49530
rect 35190 49478 35242 49530
rect 65654 49478 65706 49530
rect 65718 49478 65770 49530
rect 65782 49478 65834 49530
rect 65846 49478 65898 49530
rect 65910 49478 65962 49530
rect 19574 48934 19626 48986
rect 19638 48934 19690 48986
rect 19702 48934 19754 48986
rect 19766 48934 19818 48986
rect 19830 48934 19882 48986
rect 50294 48934 50346 48986
rect 50358 48934 50410 48986
rect 50422 48934 50474 48986
rect 50486 48934 50538 48986
rect 50550 48934 50602 48986
rect 4214 48390 4266 48442
rect 4278 48390 4330 48442
rect 4342 48390 4394 48442
rect 4406 48390 4458 48442
rect 4470 48390 4522 48442
rect 34934 48390 34986 48442
rect 34998 48390 35050 48442
rect 35062 48390 35114 48442
rect 35126 48390 35178 48442
rect 35190 48390 35242 48442
rect 65654 48390 65706 48442
rect 65718 48390 65770 48442
rect 65782 48390 65834 48442
rect 65846 48390 65898 48442
rect 65910 48390 65962 48442
rect 39856 48220 39908 48272
rect 75828 48220 75880 48272
rect 19574 47846 19626 47898
rect 19638 47846 19690 47898
rect 19702 47846 19754 47898
rect 19766 47846 19818 47898
rect 19830 47846 19882 47898
rect 50294 47846 50346 47898
rect 50358 47846 50410 47898
rect 50422 47846 50474 47898
rect 50486 47846 50538 47898
rect 50550 47846 50602 47898
rect 4214 47302 4266 47354
rect 4278 47302 4330 47354
rect 4342 47302 4394 47354
rect 4406 47302 4458 47354
rect 4470 47302 4522 47354
rect 34934 47302 34986 47354
rect 34998 47302 35050 47354
rect 35062 47302 35114 47354
rect 35126 47302 35178 47354
rect 35190 47302 35242 47354
rect 65654 47302 65706 47354
rect 65718 47302 65770 47354
rect 65782 47302 65834 47354
rect 65846 47302 65898 47354
rect 65910 47302 65962 47354
rect 1584 47175 1636 47184
rect 1584 47141 1593 47175
rect 1593 47141 1627 47175
rect 1627 47141 1636 47175
rect 1584 47132 1636 47141
rect 2872 46996 2924 47048
rect 19574 46758 19626 46810
rect 19638 46758 19690 46810
rect 19702 46758 19754 46810
rect 19766 46758 19818 46810
rect 19830 46758 19882 46810
rect 50294 46758 50346 46810
rect 50358 46758 50410 46810
rect 50422 46758 50474 46810
rect 50486 46758 50538 46810
rect 50550 46758 50602 46810
rect 4214 46214 4266 46266
rect 4278 46214 4330 46266
rect 4342 46214 4394 46266
rect 4406 46214 4458 46266
rect 4470 46214 4522 46266
rect 34934 46214 34986 46266
rect 34998 46214 35050 46266
rect 35062 46214 35114 46266
rect 35126 46214 35178 46266
rect 35190 46214 35242 46266
rect 65654 46214 65706 46266
rect 65718 46214 65770 46266
rect 65782 46214 65834 46266
rect 65846 46214 65898 46266
rect 65910 46214 65962 46266
rect 19574 45670 19626 45722
rect 19638 45670 19690 45722
rect 19702 45670 19754 45722
rect 19766 45670 19818 45722
rect 19830 45670 19882 45722
rect 50294 45670 50346 45722
rect 50358 45670 50410 45722
rect 50422 45670 50474 45722
rect 50486 45670 50538 45722
rect 50550 45670 50602 45722
rect 4214 45126 4266 45178
rect 4278 45126 4330 45178
rect 4342 45126 4394 45178
rect 4406 45126 4458 45178
rect 4470 45126 4522 45178
rect 34934 45126 34986 45178
rect 34998 45126 35050 45178
rect 35062 45126 35114 45178
rect 35126 45126 35178 45178
rect 35190 45126 35242 45178
rect 65654 45126 65706 45178
rect 65718 45126 65770 45178
rect 65782 45126 65834 45178
rect 65846 45126 65898 45178
rect 65910 45126 65962 45178
rect 19574 44582 19626 44634
rect 19638 44582 19690 44634
rect 19702 44582 19754 44634
rect 19766 44582 19818 44634
rect 19830 44582 19882 44634
rect 50294 44582 50346 44634
rect 50358 44582 50410 44634
rect 50422 44582 50474 44634
rect 50486 44582 50538 44634
rect 50550 44582 50602 44634
rect 4214 44038 4266 44090
rect 4278 44038 4330 44090
rect 4342 44038 4394 44090
rect 4406 44038 4458 44090
rect 4470 44038 4522 44090
rect 34934 44038 34986 44090
rect 34998 44038 35050 44090
rect 35062 44038 35114 44090
rect 35126 44038 35178 44090
rect 35190 44038 35242 44090
rect 65654 44038 65706 44090
rect 65718 44038 65770 44090
rect 65782 44038 65834 44090
rect 65846 44038 65898 44090
rect 65910 44038 65962 44090
rect 76564 43732 76616 43784
rect 78036 43639 78088 43648
rect 78036 43605 78045 43639
rect 78045 43605 78079 43639
rect 78079 43605 78088 43639
rect 78036 43596 78088 43605
rect 19574 43494 19626 43546
rect 19638 43494 19690 43546
rect 19702 43494 19754 43546
rect 19766 43494 19818 43546
rect 19830 43494 19882 43546
rect 50294 43494 50346 43546
rect 50358 43494 50410 43546
rect 50422 43494 50474 43546
rect 50486 43494 50538 43546
rect 50550 43494 50602 43546
rect 1860 43299 1912 43308
rect 1860 43265 1869 43299
rect 1869 43265 1903 43299
rect 1903 43265 1912 43299
rect 1860 43256 1912 43265
rect 39580 43052 39632 43104
rect 4214 42950 4266 43002
rect 4278 42950 4330 43002
rect 4342 42950 4394 43002
rect 4406 42950 4458 43002
rect 4470 42950 4522 43002
rect 34934 42950 34986 43002
rect 34998 42950 35050 43002
rect 35062 42950 35114 43002
rect 35126 42950 35178 43002
rect 35190 42950 35242 43002
rect 65654 42950 65706 43002
rect 65718 42950 65770 43002
rect 65782 42950 65834 43002
rect 65846 42950 65898 43002
rect 65910 42950 65962 43002
rect 77760 42755 77812 42764
rect 77760 42721 77769 42755
rect 77769 42721 77803 42755
rect 77803 42721 77812 42755
rect 77760 42712 77812 42721
rect 77576 42619 77628 42628
rect 77576 42585 77585 42619
rect 77585 42585 77619 42619
rect 77619 42585 77628 42619
rect 77576 42576 77628 42585
rect 19574 42406 19626 42458
rect 19638 42406 19690 42458
rect 19702 42406 19754 42458
rect 19766 42406 19818 42458
rect 19830 42406 19882 42458
rect 50294 42406 50346 42458
rect 50358 42406 50410 42458
rect 50422 42406 50474 42458
rect 50486 42406 50538 42458
rect 50550 42406 50602 42458
rect 4214 41862 4266 41914
rect 4278 41862 4330 41914
rect 4342 41862 4394 41914
rect 4406 41862 4458 41914
rect 4470 41862 4522 41914
rect 34934 41862 34986 41914
rect 34998 41862 35050 41914
rect 35062 41862 35114 41914
rect 35126 41862 35178 41914
rect 35190 41862 35242 41914
rect 65654 41862 65706 41914
rect 65718 41862 65770 41914
rect 65782 41862 65834 41914
rect 65846 41862 65898 41914
rect 65910 41862 65962 41914
rect 19574 41318 19626 41370
rect 19638 41318 19690 41370
rect 19702 41318 19754 41370
rect 19766 41318 19818 41370
rect 19830 41318 19882 41370
rect 50294 41318 50346 41370
rect 50358 41318 50410 41370
rect 50422 41318 50474 41370
rect 50486 41318 50538 41370
rect 50550 41318 50602 41370
rect 4214 40774 4266 40826
rect 4278 40774 4330 40826
rect 4342 40774 4394 40826
rect 4406 40774 4458 40826
rect 4470 40774 4522 40826
rect 34934 40774 34986 40826
rect 34998 40774 35050 40826
rect 35062 40774 35114 40826
rect 35126 40774 35178 40826
rect 35190 40774 35242 40826
rect 65654 40774 65706 40826
rect 65718 40774 65770 40826
rect 65782 40774 65834 40826
rect 65846 40774 65898 40826
rect 65910 40774 65962 40826
rect 77484 40468 77536 40520
rect 78036 40375 78088 40384
rect 78036 40341 78045 40375
rect 78045 40341 78079 40375
rect 78079 40341 78088 40375
rect 78036 40332 78088 40341
rect 19574 40230 19626 40282
rect 19638 40230 19690 40282
rect 19702 40230 19754 40282
rect 19766 40230 19818 40282
rect 19830 40230 19882 40282
rect 50294 40230 50346 40282
rect 50358 40230 50410 40282
rect 50422 40230 50474 40282
rect 50486 40230 50538 40282
rect 50550 40230 50602 40282
rect 77484 40171 77536 40180
rect 77484 40137 77493 40171
rect 77493 40137 77527 40171
rect 77527 40137 77536 40171
rect 77484 40128 77536 40137
rect 77576 40060 77628 40112
rect 4214 39686 4266 39738
rect 4278 39686 4330 39738
rect 4342 39686 4394 39738
rect 4406 39686 4458 39738
rect 4470 39686 4522 39738
rect 34934 39686 34986 39738
rect 34998 39686 35050 39738
rect 35062 39686 35114 39738
rect 35126 39686 35178 39738
rect 35190 39686 35242 39738
rect 65654 39686 65706 39738
rect 65718 39686 65770 39738
rect 65782 39686 65834 39738
rect 65846 39686 65898 39738
rect 65910 39686 65962 39738
rect 19574 39142 19626 39194
rect 19638 39142 19690 39194
rect 19702 39142 19754 39194
rect 19766 39142 19818 39194
rect 19830 39142 19882 39194
rect 50294 39142 50346 39194
rect 50358 39142 50410 39194
rect 50422 39142 50474 39194
rect 50486 39142 50538 39194
rect 50550 39142 50602 39194
rect 1860 38947 1912 38956
rect 1860 38913 1869 38947
rect 1869 38913 1903 38947
rect 1903 38913 1912 38947
rect 1860 38904 1912 38913
rect 38844 38700 38896 38752
rect 4214 38598 4266 38650
rect 4278 38598 4330 38650
rect 4342 38598 4394 38650
rect 4406 38598 4458 38650
rect 4470 38598 4522 38650
rect 34934 38598 34986 38650
rect 34998 38598 35050 38650
rect 35062 38598 35114 38650
rect 35126 38598 35178 38650
rect 35190 38598 35242 38650
rect 65654 38598 65706 38650
rect 65718 38598 65770 38650
rect 65782 38598 65834 38650
rect 65846 38598 65898 38650
rect 65910 38598 65962 38650
rect 19574 38054 19626 38106
rect 19638 38054 19690 38106
rect 19702 38054 19754 38106
rect 19766 38054 19818 38106
rect 19830 38054 19882 38106
rect 50294 38054 50346 38106
rect 50358 38054 50410 38106
rect 50422 38054 50474 38106
rect 50486 38054 50538 38106
rect 50550 38054 50602 38106
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 34934 37510 34986 37562
rect 34998 37510 35050 37562
rect 35062 37510 35114 37562
rect 35126 37510 35178 37562
rect 35190 37510 35242 37562
rect 65654 37510 65706 37562
rect 65718 37510 65770 37562
rect 65782 37510 65834 37562
rect 65846 37510 65898 37562
rect 65910 37510 65962 37562
rect 19574 36966 19626 37018
rect 19638 36966 19690 37018
rect 19702 36966 19754 37018
rect 19766 36966 19818 37018
rect 19830 36966 19882 37018
rect 50294 36966 50346 37018
rect 50358 36966 50410 37018
rect 50422 36966 50474 37018
rect 50486 36966 50538 37018
rect 50550 36966 50602 37018
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 65654 36422 65706 36474
rect 65718 36422 65770 36474
rect 65782 36422 65834 36474
rect 65846 36422 65898 36474
rect 65910 36422 65962 36474
rect 77852 36159 77904 36168
rect 77852 36125 77861 36159
rect 77861 36125 77895 36159
rect 77895 36125 77904 36159
rect 77852 36116 77904 36125
rect 78036 36023 78088 36032
rect 78036 35989 78045 36023
rect 78045 35989 78079 36023
rect 78079 35989 78088 36023
rect 78036 35980 78088 35989
rect 19574 35878 19626 35930
rect 19638 35878 19690 35930
rect 19702 35878 19754 35930
rect 19766 35878 19818 35930
rect 19830 35878 19882 35930
rect 50294 35878 50346 35930
rect 50358 35878 50410 35930
rect 50422 35878 50474 35930
rect 50486 35878 50538 35930
rect 50550 35878 50602 35930
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 65654 35334 65706 35386
rect 65718 35334 65770 35386
rect 65782 35334 65834 35386
rect 65846 35334 65898 35386
rect 65910 35334 65962 35386
rect 1492 35028 1544 35080
rect 1584 34935 1636 34944
rect 1584 34901 1593 34935
rect 1593 34901 1627 34935
rect 1627 34901 1636 34935
rect 1584 34892 1636 34901
rect 19574 34790 19626 34842
rect 19638 34790 19690 34842
rect 19702 34790 19754 34842
rect 19766 34790 19818 34842
rect 19830 34790 19882 34842
rect 50294 34790 50346 34842
rect 50358 34790 50410 34842
rect 50422 34790 50474 34842
rect 50486 34790 50538 34842
rect 50550 34790 50602 34842
rect 76564 34620 76616 34672
rect 66628 34552 66680 34604
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 65654 34246 65706 34298
rect 65718 34246 65770 34298
rect 65782 34246 65834 34298
rect 65846 34246 65898 34298
rect 65910 34246 65962 34298
rect 19574 33702 19626 33754
rect 19638 33702 19690 33754
rect 19702 33702 19754 33754
rect 19766 33702 19818 33754
rect 19830 33702 19882 33754
rect 50294 33702 50346 33754
rect 50358 33702 50410 33754
rect 50422 33702 50474 33754
rect 50486 33702 50538 33754
rect 50550 33702 50602 33754
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 65654 33158 65706 33210
rect 65718 33158 65770 33210
rect 65782 33158 65834 33210
rect 65846 33158 65898 33210
rect 65910 33158 65962 33210
rect 77852 33099 77904 33108
rect 77852 33065 77861 33099
rect 77861 33065 77895 33099
rect 77895 33065 77904 33099
rect 77852 33056 77904 33065
rect 78036 32895 78088 32904
rect 78036 32861 78045 32895
rect 78045 32861 78079 32895
rect 78079 32861 78088 32895
rect 78036 32852 78088 32861
rect 19574 32614 19626 32666
rect 19638 32614 19690 32666
rect 19702 32614 19754 32666
rect 19766 32614 19818 32666
rect 19830 32614 19882 32666
rect 50294 32614 50346 32666
rect 50358 32614 50410 32666
rect 50422 32614 50474 32666
rect 50486 32614 50538 32666
rect 50550 32614 50602 32666
rect 77760 32376 77812 32428
rect 77852 32215 77904 32224
rect 77852 32181 77861 32215
rect 77861 32181 77895 32215
rect 77895 32181 77904 32215
rect 77852 32172 77904 32181
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 65654 32070 65706 32122
rect 65718 32070 65770 32122
rect 65782 32070 65834 32122
rect 65846 32070 65898 32122
rect 65910 32070 65962 32122
rect 40776 31832 40828 31884
rect 1400 31807 1452 31816
rect 1400 31773 1409 31807
rect 1409 31773 1443 31807
rect 1443 31773 1452 31807
rect 1400 31764 1452 31773
rect 19574 31526 19626 31578
rect 19638 31526 19690 31578
rect 19702 31526 19754 31578
rect 19766 31526 19818 31578
rect 19830 31526 19882 31578
rect 50294 31526 50346 31578
rect 50358 31526 50410 31578
rect 50422 31526 50474 31578
rect 50486 31526 50538 31578
rect 50550 31526 50602 31578
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 65654 30982 65706 31034
rect 65718 30982 65770 31034
rect 65782 30982 65834 31034
rect 65846 30982 65898 31034
rect 65910 30982 65962 31034
rect 19574 30438 19626 30490
rect 19638 30438 19690 30490
rect 19702 30438 19754 30490
rect 19766 30438 19818 30490
rect 19830 30438 19882 30490
rect 50294 30438 50346 30490
rect 50358 30438 50410 30490
rect 50422 30438 50474 30490
rect 50486 30438 50538 30490
rect 50550 30438 50602 30490
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 65654 29894 65706 29946
rect 65718 29894 65770 29946
rect 65782 29894 65834 29946
rect 65846 29894 65898 29946
rect 65910 29894 65962 29946
rect 19574 29350 19626 29402
rect 19638 29350 19690 29402
rect 19702 29350 19754 29402
rect 19766 29350 19818 29402
rect 19830 29350 19882 29402
rect 50294 29350 50346 29402
rect 50358 29350 50410 29402
rect 50422 29350 50474 29402
rect 50486 29350 50538 29402
rect 50550 29350 50602 29402
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 65654 28806 65706 28858
rect 65718 28806 65770 28858
rect 65782 28806 65834 28858
rect 65846 28806 65898 28858
rect 65910 28806 65962 28858
rect 19574 28262 19626 28314
rect 19638 28262 19690 28314
rect 19702 28262 19754 28314
rect 19766 28262 19818 28314
rect 19830 28262 19882 28314
rect 50294 28262 50346 28314
rect 50358 28262 50410 28314
rect 50422 28262 50474 28314
rect 50486 28262 50538 28314
rect 50550 28262 50602 28314
rect 78036 28160 78088 28212
rect 77944 28067 77996 28076
rect 77944 28033 77953 28067
rect 77953 28033 77987 28067
rect 77987 28033 77996 28067
rect 77944 28024 77996 28033
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 65654 27718 65706 27770
rect 65718 27718 65770 27770
rect 65782 27718 65834 27770
rect 65846 27718 65898 27770
rect 65910 27718 65962 27770
rect 1400 27455 1452 27464
rect 1400 27421 1409 27455
rect 1409 27421 1443 27455
rect 1443 27421 1452 27455
rect 1400 27412 1452 27421
rect 39672 27344 39724 27396
rect 19574 27174 19626 27226
rect 19638 27174 19690 27226
rect 19702 27174 19754 27226
rect 19766 27174 19818 27226
rect 19830 27174 19882 27226
rect 50294 27174 50346 27226
rect 50358 27174 50410 27226
rect 50422 27174 50474 27226
rect 50486 27174 50538 27226
rect 50550 27174 50602 27226
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 65654 26630 65706 26682
rect 65718 26630 65770 26682
rect 65782 26630 65834 26682
rect 65846 26630 65898 26682
rect 65910 26630 65962 26682
rect 19574 26086 19626 26138
rect 19638 26086 19690 26138
rect 19702 26086 19754 26138
rect 19766 26086 19818 26138
rect 19830 26086 19882 26138
rect 50294 26086 50346 26138
rect 50358 26086 50410 26138
rect 50422 26086 50474 26138
rect 50486 26086 50538 26138
rect 50550 26086 50602 26138
rect 77852 25848 77904 25900
rect 39580 25644 39632 25696
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 65654 25542 65706 25594
rect 65718 25542 65770 25594
rect 65782 25542 65834 25594
rect 65846 25542 65898 25594
rect 65910 25542 65962 25594
rect 1768 25440 1820 25492
rect 39580 25440 39632 25492
rect 19574 24998 19626 25050
rect 19638 24998 19690 25050
rect 19702 24998 19754 25050
rect 19766 24998 19818 25050
rect 19830 24998 19882 25050
rect 50294 24998 50346 25050
rect 50358 24998 50410 25050
rect 50422 24998 50474 25050
rect 50486 24998 50538 25050
rect 50550 24998 50602 25050
rect 39120 24556 39172 24608
rect 77852 24599 77904 24608
rect 77852 24565 77861 24599
rect 77861 24565 77895 24599
rect 77895 24565 77904 24599
rect 77852 24556 77904 24565
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 65654 24454 65706 24506
rect 65718 24454 65770 24506
rect 65782 24454 65834 24506
rect 65846 24454 65898 24506
rect 65910 24454 65962 24506
rect 19574 23910 19626 23962
rect 19638 23910 19690 23962
rect 19702 23910 19754 23962
rect 19766 23910 19818 23962
rect 19830 23910 19882 23962
rect 50294 23910 50346 23962
rect 50358 23910 50410 23962
rect 50422 23910 50474 23962
rect 50486 23910 50538 23962
rect 50550 23910 50602 23962
rect 1400 23715 1452 23724
rect 1400 23681 1409 23715
rect 1409 23681 1443 23715
rect 1443 23681 1452 23715
rect 1400 23672 1452 23681
rect 38936 23604 38988 23656
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 65654 23366 65706 23418
rect 65718 23366 65770 23418
rect 65782 23366 65834 23418
rect 65846 23366 65898 23418
rect 65910 23366 65962 23418
rect 19574 22822 19626 22874
rect 19638 22822 19690 22874
rect 19702 22822 19754 22874
rect 19766 22822 19818 22874
rect 19830 22822 19882 22874
rect 50294 22822 50346 22874
rect 50358 22822 50410 22874
rect 50422 22822 50474 22874
rect 50486 22822 50538 22874
rect 50550 22822 50602 22874
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 65654 22278 65706 22330
rect 65718 22278 65770 22330
rect 65782 22278 65834 22330
rect 65846 22278 65898 22330
rect 65910 22278 65962 22330
rect 19574 21734 19626 21786
rect 19638 21734 19690 21786
rect 19702 21734 19754 21786
rect 19766 21734 19818 21786
rect 19830 21734 19882 21786
rect 50294 21734 50346 21786
rect 50358 21734 50410 21786
rect 50422 21734 50474 21786
rect 50486 21734 50538 21786
rect 50550 21734 50602 21786
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 65654 21190 65706 21242
rect 65718 21190 65770 21242
rect 65782 21190 65834 21242
rect 65846 21190 65898 21242
rect 65910 21190 65962 21242
rect 77760 20884 77812 20936
rect 78036 20791 78088 20800
rect 78036 20757 78045 20791
rect 78045 20757 78079 20791
rect 78079 20757 78088 20791
rect 78036 20748 78088 20757
rect 19574 20646 19626 20698
rect 19638 20646 19690 20698
rect 19702 20646 19754 20698
rect 19766 20646 19818 20698
rect 19830 20646 19882 20698
rect 50294 20646 50346 20698
rect 50358 20646 50410 20698
rect 50422 20646 50474 20698
rect 50486 20646 50538 20698
rect 50550 20646 50602 20698
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 65654 20102 65706 20154
rect 65718 20102 65770 20154
rect 65782 20102 65834 20154
rect 65846 20102 65898 20154
rect 65910 20102 65962 20154
rect 19574 19558 19626 19610
rect 19638 19558 19690 19610
rect 19702 19558 19754 19610
rect 19766 19558 19818 19610
rect 19830 19558 19882 19610
rect 50294 19558 50346 19610
rect 50358 19558 50410 19610
rect 50422 19558 50474 19610
rect 50486 19558 50538 19610
rect 50550 19558 50602 19610
rect 1492 19320 1544 19372
rect 1584 19159 1636 19168
rect 1584 19125 1593 19159
rect 1593 19125 1627 19159
rect 1627 19125 1636 19159
rect 1584 19116 1636 19125
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 65654 19014 65706 19066
rect 65718 19014 65770 19066
rect 65782 19014 65834 19066
rect 65846 19014 65898 19066
rect 65910 19014 65962 19066
rect 19574 18470 19626 18522
rect 19638 18470 19690 18522
rect 19702 18470 19754 18522
rect 19766 18470 19818 18522
rect 19830 18470 19882 18522
rect 50294 18470 50346 18522
rect 50358 18470 50410 18522
rect 50422 18470 50474 18522
rect 50486 18470 50538 18522
rect 50550 18470 50602 18522
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 65654 17926 65706 17978
rect 65718 17926 65770 17978
rect 65782 17926 65834 17978
rect 65846 17926 65898 17978
rect 65910 17926 65962 17978
rect 19574 17382 19626 17434
rect 19638 17382 19690 17434
rect 19702 17382 19754 17434
rect 19766 17382 19818 17434
rect 19830 17382 19882 17434
rect 50294 17382 50346 17434
rect 50358 17382 50410 17434
rect 50422 17382 50474 17434
rect 50486 17382 50538 17434
rect 50550 17382 50602 17434
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 65654 16838 65706 16890
rect 65718 16838 65770 16890
rect 65782 16838 65834 16890
rect 65846 16838 65898 16890
rect 65910 16838 65962 16890
rect 63040 16532 63092 16584
rect 78036 16439 78088 16448
rect 78036 16405 78045 16439
rect 78045 16405 78079 16439
rect 78079 16405 78088 16439
rect 78036 16396 78088 16405
rect 19574 16294 19626 16346
rect 19638 16294 19690 16346
rect 19702 16294 19754 16346
rect 19766 16294 19818 16346
rect 19830 16294 19882 16346
rect 50294 16294 50346 16346
rect 50358 16294 50410 16346
rect 50422 16294 50474 16346
rect 50486 16294 50538 16346
rect 50550 16294 50602 16346
rect 1768 16192 1820 16244
rect 1492 15895 1544 15904
rect 1492 15861 1501 15895
rect 1501 15861 1535 15895
rect 1535 15861 1544 15895
rect 1492 15852 1544 15861
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 65654 15750 65706 15802
rect 65718 15750 65770 15802
rect 65782 15750 65834 15802
rect 65846 15750 65898 15802
rect 65910 15750 65962 15802
rect 19574 15206 19626 15258
rect 19638 15206 19690 15258
rect 19702 15206 19754 15258
rect 19766 15206 19818 15258
rect 19830 15206 19882 15258
rect 50294 15206 50346 15258
rect 50358 15206 50410 15258
rect 50422 15206 50474 15258
rect 50486 15206 50538 15258
rect 50550 15206 50602 15258
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 65654 14662 65706 14714
rect 65718 14662 65770 14714
rect 65782 14662 65834 14714
rect 65846 14662 65898 14714
rect 65910 14662 65962 14714
rect 19574 14118 19626 14170
rect 19638 14118 19690 14170
rect 19702 14118 19754 14170
rect 19766 14118 19818 14170
rect 19830 14118 19882 14170
rect 50294 14118 50346 14170
rect 50358 14118 50410 14170
rect 50422 14118 50474 14170
rect 50486 14118 50538 14170
rect 50550 14118 50602 14170
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 65654 13574 65706 13626
rect 65718 13574 65770 13626
rect 65782 13574 65834 13626
rect 65846 13574 65898 13626
rect 65910 13574 65962 13626
rect 2872 13515 2924 13524
rect 2872 13481 2881 13515
rect 2881 13481 2915 13515
rect 2915 13481 2924 13515
rect 2872 13472 2924 13481
rect 2412 13268 2464 13320
rect 19574 13030 19626 13082
rect 19638 13030 19690 13082
rect 19702 13030 19754 13082
rect 19766 13030 19818 13082
rect 19830 13030 19882 13082
rect 50294 13030 50346 13082
rect 50358 13030 50410 13082
rect 50422 13030 50474 13082
rect 50486 13030 50538 13082
rect 50550 13030 50602 13082
rect 77668 12860 77720 12912
rect 77208 12792 77260 12844
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 65654 12486 65706 12538
rect 65718 12486 65770 12538
rect 65782 12486 65834 12538
rect 65846 12486 65898 12538
rect 65910 12486 65962 12538
rect 18328 12112 18380 12164
rect 77760 12044 77812 12096
rect 19574 11942 19626 11994
rect 19638 11942 19690 11994
rect 19702 11942 19754 11994
rect 19766 11942 19818 11994
rect 19830 11942 19882 11994
rect 50294 11942 50346 11994
rect 50358 11942 50410 11994
rect 50422 11942 50474 11994
rect 50486 11942 50538 11994
rect 50550 11942 50602 11994
rect 3056 11772 3108 11824
rect 1400 11747 1452 11756
rect 1400 11713 1409 11747
rect 1409 11713 1443 11747
rect 1443 11713 1452 11747
rect 1400 11704 1452 11713
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 65654 11398 65706 11450
rect 65718 11398 65770 11450
rect 65782 11398 65834 11450
rect 65846 11398 65898 11450
rect 65910 11398 65962 11450
rect 19574 10854 19626 10906
rect 19638 10854 19690 10906
rect 19702 10854 19754 10906
rect 19766 10854 19818 10906
rect 19830 10854 19882 10906
rect 50294 10854 50346 10906
rect 50358 10854 50410 10906
rect 50422 10854 50474 10906
rect 50486 10854 50538 10906
rect 50550 10854 50602 10906
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 65654 10310 65706 10362
rect 65718 10310 65770 10362
rect 65782 10310 65834 10362
rect 65846 10310 65898 10362
rect 65910 10310 65962 10362
rect 78128 10072 78180 10124
rect 77944 10004 77996 10056
rect 19574 9766 19626 9818
rect 19638 9766 19690 9818
rect 19702 9766 19754 9818
rect 19766 9766 19818 9818
rect 19830 9766 19882 9818
rect 50294 9766 50346 9818
rect 50358 9766 50410 9818
rect 50422 9766 50474 9818
rect 50486 9766 50538 9818
rect 50550 9766 50602 9818
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 65654 9222 65706 9274
rect 65718 9222 65770 9274
rect 65782 9222 65834 9274
rect 65846 9222 65898 9274
rect 65910 9222 65962 9274
rect 40592 8780 40644 8832
rect 78036 8823 78088 8832
rect 78036 8789 78045 8823
rect 78045 8789 78079 8823
rect 78079 8789 78088 8823
rect 78036 8780 78088 8789
rect 19574 8678 19626 8730
rect 19638 8678 19690 8730
rect 19702 8678 19754 8730
rect 19766 8678 19818 8730
rect 19830 8678 19882 8730
rect 50294 8678 50346 8730
rect 50358 8678 50410 8730
rect 50422 8678 50474 8730
rect 50486 8678 50538 8730
rect 50550 8678 50602 8730
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 65654 8134 65706 8186
rect 65718 8134 65770 8186
rect 65782 8134 65834 8186
rect 65846 8134 65898 8186
rect 65910 8134 65962 8186
rect 2688 7828 2740 7880
rect 1584 7735 1636 7744
rect 1584 7701 1593 7735
rect 1593 7701 1627 7735
rect 1627 7701 1636 7735
rect 1584 7692 1636 7701
rect 19574 7590 19626 7642
rect 19638 7590 19690 7642
rect 19702 7590 19754 7642
rect 19766 7590 19818 7642
rect 19830 7590 19882 7642
rect 50294 7590 50346 7642
rect 50358 7590 50410 7642
rect 50422 7590 50474 7642
rect 50486 7590 50538 7642
rect 50550 7590 50602 7642
rect 2412 7531 2464 7540
rect 2412 7497 2421 7531
rect 2421 7497 2455 7531
rect 2455 7497 2464 7531
rect 2412 7488 2464 7497
rect 2688 7531 2740 7540
rect 2688 7497 2697 7531
rect 2697 7497 2731 7531
rect 2731 7497 2740 7531
rect 2688 7488 2740 7497
rect 29920 7352 29972 7404
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 65654 7046 65706 7098
rect 65718 7046 65770 7098
rect 65782 7046 65834 7098
rect 65846 7046 65898 7098
rect 65910 7046 65962 7098
rect 19574 6502 19626 6554
rect 19638 6502 19690 6554
rect 19702 6502 19754 6554
rect 19766 6502 19818 6554
rect 19830 6502 19882 6554
rect 50294 6502 50346 6554
rect 50358 6502 50410 6554
rect 50422 6502 50474 6554
rect 50486 6502 50538 6554
rect 50550 6502 50602 6554
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 65654 5958 65706 6010
rect 65718 5958 65770 6010
rect 65782 5958 65834 6010
rect 65846 5958 65898 6010
rect 65910 5958 65962 6010
rect 19574 5414 19626 5466
rect 19638 5414 19690 5466
rect 19702 5414 19754 5466
rect 19766 5414 19818 5466
rect 19830 5414 19882 5466
rect 50294 5414 50346 5466
rect 50358 5414 50410 5466
rect 50422 5414 50474 5466
rect 50486 5414 50538 5466
rect 50550 5414 50602 5466
rect 77668 5219 77720 5228
rect 77668 5185 77677 5219
rect 77677 5185 77711 5219
rect 77711 5185 77720 5219
rect 77668 5176 77720 5185
rect 77852 5015 77904 5024
rect 77852 4981 77861 5015
rect 77861 4981 77895 5015
rect 77895 4981 77904 5015
rect 77852 4972 77904 4981
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 65654 4870 65706 4922
rect 65718 4870 65770 4922
rect 65782 4870 65834 4922
rect 65846 4870 65898 4922
rect 65910 4870 65962 4922
rect 77668 4768 77720 4820
rect 78036 4607 78088 4616
rect 78036 4573 78045 4607
rect 78045 4573 78079 4607
rect 78079 4573 78088 4607
rect 78036 4564 78088 4573
rect 19574 4326 19626 4378
rect 19638 4326 19690 4378
rect 19702 4326 19754 4378
rect 19766 4326 19818 4378
rect 19830 4326 19882 4378
rect 50294 4326 50346 4378
rect 50358 4326 50410 4378
rect 50422 4326 50474 4378
rect 50486 4326 50538 4378
rect 50550 4326 50602 4378
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 65654 3782 65706 3834
rect 65718 3782 65770 3834
rect 65782 3782 65834 3834
rect 65846 3782 65898 3834
rect 65910 3782 65962 3834
rect 1676 3587 1728 3596
rect 1676 3553 1685 3587
rect 1685 3553 1719 3587
rect 1719 3553 1728 3587
rect 1676 3544 1728 3553
rect 1400 3519 1452 3528
rect 1400 3485 1409 3519
rect 1409 3485 1443 3519
rect 1443 3485 1452 3519
rect 1400 3476 1452 3485
rect 12440 3476 12492 3528
rect 40960 3519 41012 3528
rect 40960 3485 40969 3519
rect 40969 3485 41003 3519
rect 41003 3485 41012 3519
rect 40960 3476 41012 3485
rect 43904 3476 43956 3528
rect 57980 3408 58032 3460
rect 16212 3340 16264 3392
rect 40408 3383 40460 3392
rect 40408 3349 40417 3383
rect 40417 3349 40451 3383
rect 40451 3349 40460 3383
rect 40408 3340 40460 3349
rect 41144 3383 41196 3392
rect 41144 3349 41153 3383
rect 41153 3349 41187 3383
rect 41187 3349 41196 3383
rect 41144 3340 41196 3349
rect 41696 3383 41748 3392
rect 41696 3349 41705 3383
rect 41705 3349 41739 3383
rect 41739 3349 41748 3383
rect 41696 3340 41748 3349
rect 19574 3238 19626 3290
rect 19638 3238 19690 3290
rect 19702 3238 19754 3290
rect 19766 3238 19818 3290
rect 19830 3238 19882 3290
rect 50294 3238 50346 3290
rect 50358 3238 50410 3290
rect 50422 3238 50474 3290
rect 50486 3238 50538 3290
rect 50550 3238 50602 3290
rect 11520 3136 11572 3188
rect 40408 3136 40460 3188
rect 77668 3000 77720 3052
rect 41236 2932 41288 2984
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 65654 2694 65706 2746
rect 65718 2694 65770 2746
rect 65782 2694 65834 2746
rect 65846 2694 65898 2746
rect 65910 2694 65962 2746
rect 18328 2635 18380 2644
rect 18328 2601 18337 2635
rect 18337 2601 18371 2635
rect 18371 2601 18380 2635
rect 18328 2592 18380 2601
rect 29920 2635 29972 2644
rect 29920 2601 29929 2635
rect 29929 2601 29963 2635
rect 29963 2601 29972 2635
rect 29920 2592 29972 2601
rect 33140 2635 33192 2644
rect 33140 2601 33149 2635
rect 33149 2601 33183 2635
rect 33183 2601 33192 2635
rect 33140 2592 33192 2601
rect 12440 2524 12492 2576
rect 40960 2592 41012 2644
rect 43904 2592 43956 2644
rect 41052 2524 41104 2576
rect 55772 2592 55824 2644
rect 66628 2635 66680 2644
rect 66628 2601 66637 2635
rect 66637 2601 66671 2635
rect 66671 2601 66680 2635
rect 66628 2592 66680 2601
rect 50620 2524 50672 2576
rect 4620 2456 4672 2508
rect 19984 2456 20036 2508
rect 20 2388 72 2440
rect 3240 2388 3292 2440
rect 7104 2388 7156 2440
rect 11520 2431 11572 2440
rect 11520 2397 11529 2431
rect 11529 2397 11563 2431
rect 11563 2397 11572 2431
rect 11520 2388 11572 2397
rect 16212 2388 16264 2440
rect 41144 2456 41196 2508
rect 29644 2388 29696 2440
rect 35348 2388 35400 2440
rect 41696 2388 41748 2440
rect 44456 2388 44508 2440
rect 47676 2388 47728 2440
rect 51540 2388 51592 2440
rect 55404 2388 55456 2440
rect 55772 2431 55824 2440
rect 55772 2397 55781 2431
rect 55781 2397 55815 2431
rect 55815 2397 55824 2431
rect 55772 2388 55824 2397
rect 59268 2388 59320 2440
rect 7840 2363 7892 2372
rect 7840 2329 7849 2363
rect 7849 2329 7883 2363
rect 7883 2329 7892 2363
rect 7840 2320 7892 2329
rect 14832 2320 14884 2372
rect 18052 2320 18104 2372
rect 32864 2320 32916 2372
rect 39764 2320 39816 2372
rect 51908 2363 51960 2372
rect 51908 2329 51917 2363
rect 51917 2329 51951 2363
rect 51951 2329 51960 2363
rect 51908 2320 51960 2329
rect 57980 2320 58032 2372
rect 62488 2388 62540 2440
rect 66352 2388 66404 2440
rect 70216 2388 70268 2440
rect 78036 2456 78088 2508
rect 77300 2388 77352 2440
rect 63868 2363 63920 2372
rect 63868 2329 63877 2363
rect 63877 2329 63911 2363
rect 63911 2329 63920 2363
rect 63868 2320 63920 2329
rect 10968 2252 11020 2304
rect 21916 2252 21968 2304
rect 25780 2252 25832 2304
rect 36728 2252 36780 2304
rect 40592 2252 40644 2304
rect 40960 2252 41012 2304
rect 50620 2252 50672 2304
rect 74080 2252 74132 2304
rect 19574 2150 19626 2202
rect 19638 2150 19690 2202
rect 19702 2150 19754 2202
rect 19766 2150 19818 2202
rect 19830 2150 19882 2202
rect 50294 2150 50346 2202
rect 50358 2150 50410 2202
rect 50422 2150 50474 2202
rect 50486 2150 50538 2202
rect 50550 2150 50602 2202
rect 2964 1980 3016 2032
rect 63868 1980 63920 2032
rect 39948 1912 40000 1964
rect 51908 1912 51960 1964
rect 7840 1844 7892 1896
rect 77576 1844 77628 1896
<< metal2 >>
rect 662 119200 718 120000
rect 4526 119354 4582 120000
rect 7746 119354 7802 120000
rect 11610 119354 11666 120000
rect 15474 119354 15530 120000
rect 4526 119326 4660 119354
rect 4526 119200 4582 119326
rect 676 117298 704 119200
rect 4632 117366 4660 119326
rect 7746 119326 8064 119354
rect 7746 119200 7802 119326
rect 4620 117360 4672 117366
rect 4620 117302 4672 117308
rect 664 117292 716 117298
rect 664 117234 716 117240
rect 7840 117292 7892 117298
rect 7840 117234 7892 117240
rect 2320 117088 2372 117094
rect 1858 117056 1914 117065
rect 2320 117030 2372 117036
rect 1858 116991 1914 117000
rect 1872 116686 1900 116991
rect 1860 116680 1912 116686
rect 1860 116622 1912 116628
rect 2228 116612 2280 116618
rect 2228 116554 2280 116560
rect 1400 113416 1452 113422
rect 1400 113358 1452 113364
rect 1412 113174 1440 113358
rect 1584 113280 1636 113286
rect 1584 113222 1636 113228
rect 1412 113146 1532 113174
rect 1400 105800 1452 105806
rect 1400 105742 1452 105748
rect 1412 105505 1440 105742
rect 1398 105496 1454 105505
rect 1398 105431 1454 105440
rect 1400 101448 1452 101454
rect 1398 101416 1400 101425
rect 1452 101416 1454 101425
rect 1398 101351 1454 101360
rect 1400 97708 1452 97714
rect 1400 97650 1452 97656
rect 1412 97345 1440 97650
rect 1398 97336 1454 97345
rect 1398 97271 1454 97280
rect 1504 95878 1532 113146
rect 1596 112985 1624 113222
rect 1582 112976 1638 112985
rect 1582 112911 1638 112920
rect 1860 109676 1912 109682
rect 1860 109618 1912 109624
rect 1872 109585 1900 109618
rect 1858 109576 1914 109585
rect 1858 109511 1914 109520
rect 1860 105732 1912 105738
rect 1860 105674 1912 105680
rect 1676 97640 1728 97646
rect 1676 97582 1728 97588
rect 1492 95872 1544 95878
rect 1492 95814 1544 95820
rect 1584 94240 1636 94246
rect 1584 94182 1636 94188
rect 1596 93945 1624 94182
rect 1582 93936 1638 93945
rect 1582 93871 1638 93880
rect 1492 90092 1544 90098
rect 1492 90034 1544 90040
rect 1504 89865 1532 90034
rect 1490 89856 1546 89865
rect 1490 89791 1546 89800
rect 1584 86080 1636 86086
rect 1584 86022 1636 86028
rect 1596 85785 1624 86022
rect 1582 85776 1638 85785
rect 1582 85711 1638 85720
rect 1400 81864 1452 81870
rect 1400 81806 1452 81812
rect 1412 81705 1440 81806
rect 1398 81696 1454 81705
rect 1398 81631 1454 81640
rect 1584 78464 1636 78470
rect 1584 78406 1636 78412
rect 1596 78305 1624 78406
rect 1582 78296 1638 78305
rect 1582 78231 1638 78240
rect 1688 74322 1716 97582
rect 1676 74316 1728 74322
rect 1676 74258 1728 74264
rect 1492 74248 1544 74254
rect 1492 74190 1544 74196
rect 1582 74216 1638 74225
rect 1400 70508 1452 70514
rect 1400 70450 1452 70456
rect 1412 70106 1440 70450
rect 1400 70100 1452 70106
rect 1400 70042 1452 70048
rect 1400 62892 1452 62898
rect 1400 62834 1452 62840
rect 1412 59430 1440 62834
rect 1504 60586 1532 74190
rect 1582 74151 1638 74160
rect 1596 74118 1624 74151
rect 1584 74112 1636 74118
rect 1584 74054 1636 74060
rect 1676 70916 1728 70922
rect 1676 70858 1728 70864
rect 1584 70304 1636 70310
rect 1584 70246 1636 70252
rect 1596 70145 1624 70246
rect 1582 70136 1638 70145
rect 1582 70071 1638 70080
rect 1688 69902 1716 70858
rect 1676 69896 1728 69902
rect 1676 69838 1728 69844
rect 1582 66056 1638 66065
rect 1582 65991 1584 66000
rect 1636 65991 1638 66000
rect 1584 65962 1636 65968
rect 1584 62688 1636 62694
rect 1582 62656 1584 62665
rect 1636 62656 1638 62665
rect 1582 62591 1638 62600
rect 1492 60580 1544 60586
rect 1492 60522 1544 60528
rect 1492 59968 1544 59974
rect 1492 59910 1544 59916
rect 1400 59424 1452 59430
rect 1400 59366 1452 59372
rect 1400 59016 1452 59022
rect 1400 58958 1452 58964
rect 1412 58682 1440 58958
rect 1400 58676 1452 58682
rect 1400 58618 1452 58624
rect 1504 55214 1532 59910
rect 1584 58880 1636 58886
rect 1584 58822 1636 58828
rect 1596 58585 1624 58822
rect 1582 58576 1638 58585
rect 1688 58546 1716 69838
rect 1768 65408 1820 65414
rect 1768 65350 1820 65356
rect 1582 58511 1638 58520
rect 1676 58540 1728 58546
rect 1676 58482 1728 58488
rect 1780 58426 1808 65350
rect 1872 60178 1900 105674
rect 2044 86216 2096 86222
rect 2044 86158 2096 86164
rect 1952 74316 2004 74322
rect 1952 74258 2004 74264
rect 1860 60172 1912 60178
rect 1860 60114 1912 60120
rect 1964 59634 1992 74258
rect 2056 71126 2084 86158
rect 2136 81796 2188 81802
rect 2136 81738 2188 81744
rect 2044 71120 2096 71126
rect 2044 71062 2096 71068
rect 2148 60314 2176 81738
rect 2136 60308 2188 60314
rect 2136 60250 2188 60256
rect 2240 60110 2268 116554
rect 2332 66162 2360 117030
rect 4214 116988 4522 117008
rect 4214 116986 4220 116988
rect 4276 116986 4300 116988
rect 4356 116986 4380 116988
rect 4436 116986 4460 116988
rect 4516 116986 4522 116988
rect 4276 116934 4278 116986
rect 4458 116934 4460 116986
rect 4214 116932 4220 116934
rect 4276 116932 4300 116934
rect 4356 116932 4380 116934
rect 4436 116932 4460 116934
rect 4516 116932 4522 116934
rect 4214 116912 4522 116932
rect 4214 115900 4522 115920
rect 4214 115898 4220 115900
rect 4276 115898 4300 115900
rect 4356 115898 4380 115900
rect 4436 115898 4460 115900
rect 4516 115898 4522 115900
rect 4276 115846 4278 115898
rect 4458 115846 4460 115898
rect 4214 115844 4220 115846
rect 4276 115844 4300 115846
rect 4356 115844 4380 115846
rect 4436 115844 4460 115846
rect 4516 115844 4522 115846
rect 4214 115824 4522 115844
rect 4214 114812 4522 114832
rect 4214 114810 4220 114812
rect 4276 114810 4300 114812
rect 4356 114810 4380 114812
rect 4436 114810 4460 114812
rect 4516 114810 4522 114812
rect 4276 114758 4278 114810
rect 4458 114758 4460 114810
rect 4214 114756 4220 114758
rect 4276 114756 4300 114758
rect 4356 114756 4380 114758
rect 4436 114756 4460 114758
rect 4516 114756 4522 114758
rect 4214 114736 4522 114756
rect 4214 113724 4522 113744
rect 4214 113722 4220 113724
rect 4276 113722 4300 113724
rect 4356 113722 4380 113724
rect 4436 113722 4460 113724
rect 4516 113722 4522 113724
rect 4276 113670 4278 113722
rect 4458 113670 4460 113722
rect 4214 113668 4220 113670
rect 4276 113668 4300 113670
rect 4356 113668 4380 113670
rect 4436 113668 4460 113670
rect 4516 113668 4522 113670
rect 4214 113648 4522 113668
rect 4214 112636 4522 112656
rect 4214 112634 4220 112636
rect 4276 112634 4300 112636
rect 4356 112634 4380 112636
rect 4436 112634 4460 112636
rect 4516 112634 4522 112636
rect 4276 112582 4278 112634
rect 4458 112582 4460 112634
rect 4214 112580 4220 112582
rect 4276 112580 4300 112582
rect 4356 112580 4380 112582
rect 4436 112580 4460 112582
rect 4516 112580 4522 112582
rect 4214 112560 4522 112580
rect 4214 111548 4522 111568
rect 4214 111546 4220 111548
rect 4276 111546 4300 111548
rect 4356 111546 4380 111548
rect 4436 111546 4460 111548
rect 4516 111546 4522 111548
rect 4276 111494 4278 111546
rect 4458 111494 4460 111546
rect 4214 111492 4220 111494
rect 4276 111492 4300 111494
rect 4356 111492 4380 111494
rect 4436 111492 4460 111494
rect 4516 111492 4522 111494
rect 4214 111472 4522 111492
rect 4214 110460 4522 110480
rect 4214 110458 4220 110460
rect 4276 110458 4300 110460
rect 4356 110458 4380 110460
rect 4436 110458 4460 110460
rect 4516 110458 4522 110460
rect 4276 110406 4278 110458
rect 4458 110406 4460 110458
rect 4214 110404 4220 110406
rect 4276 110404 4300 110406
rect 4356 110404 4380 110406
rect 4436 110404 4460 110406
rect 4516 110404 4522 110406
rect 4214 110384 4522 110404
rect 4214 109372 4522 109392
rect 4214 109370 4220 109372
rect 4276 109370 4300 109372
rect 4356 109370 4380 109372
rect 4436 109370 4460 109372
rect 4516 109370 4522 109372
rect 4276 109318 4278 109370
rect 4458 109318 4460 109370
rect 4214 109316 4220 109318
rect 4276 109316 4300 109318
rect 4356 109316 4380 109318
rect 4436 109316 4460 109318
rect 4516 109316 4522 109318
rect 4214 109296 4522 109316
rect 4214 108284 4522 108304
rect 4214 108282 4220 108284
rect 4276 108282 4300 108284
rect 4356 108282 4380 108284
rect 4436 108282 4460 108284
rect 4516 108282 4522 108284
rect 4276 108230 4278 108282
rect 4458 108230 4460 108282
rect 4214 108228 4220 108230
rect 4276 108228 4300 108230
rect 4356 108228 4380 108230
rect 4436 108228 4460 108230
rect 4516 108228 4522 108230
rect 4214 108208 4522 108228
rect 4214 107196 4522 107216
rect 4214 107194 4220 107196
rect 4276 107194 4300 107196
rect 4356 107194 4380 107196
rect 4436 107194 4460 107196
rect 4516 107194 4522 107196
rect 4276 107142 4278 107194
rect 4458 107142 4460 107194
rect 4214 107140 4220 107142
rect 4276 107140 4300 107142
rect 4356 107140 4380 107142
rect 4436 107140 4460 107142
rect 4516 107140 4522 107142
rect 4214 107120 4522 107140
rect 4214 106108 4522 106128
rect 4214 106106 4220 106108
rect 4276 106106 4300 106108
rect 4356 106106 4380 106108
rect 4436 106106 4460 106108
rect 4516 106106 4522 106108
rect 4276 106054 4278 106106
rect 4458 106054 4460 106106
rect 4214 106052 4220 106054
rect 4276 106052 4300 106054
rect 4356 106052 4380 106054
rect 4436 106052 4460 106054
rect 4516 106052 4522 106054
rect 4214 106032 4522 106052
rect 4214 105020 4522 105040
rect 4214 105018 4220 105020
rect 4276 105018 4300 105020
rect 4356 105018 4380 105020
rect 4436 105018 4460 105020
rect 4516 105018 4522 105020
rect 4276 104966 4278 105018
rect 4458 104966 4460 105018
rect 4214 104964 4220 104966
rect 4276 104964 4300 104966
rect 4356 104964 4380 104966
rect 4436 104964 4460 104966
rect 4516 104964 4522 104966
rect 4214 104944 4522 104964
rect 4214 103932 4522 103952
rect 4214 103930 4220 103932
rect 4276 103930 4300 103932
rect 4356 103930 4380 103932
rect 4436 103930 4460 103932
rect 4516 103930 4522 103932
rect 4276 103878 4278 103930
rect 4458 103878 4460 103930
rect 4214 103876 4220 103878
rect 4276 103876 4300 103878
rect 4356 103876 4380 103878
rect 4436 103876 4460 103878
rect 4516 103876 4522 103878
rect 4214 103856 4522 103876
rect 4214 102844 4522 102864
rect 4214 102842 4220 102844
rect 4276 102842 4300 102844
rect 4356 102842 4380 102844
rect 4436 102842 4460 102844
rect 4516 102842 4522 102844
rect 4276 102790 4278 102842
rect 4458 102790 4460 102842
rect 4214 102788 4220 102790
rect 4276 102788 4300 102790
rect 4356 102788 4380 102790
rect 4436 102788 4460 102790
rect 4516 102788 4522 102790
rect 4214 102768 4522 102788
rect 4214 101756 4522 101776
rect 4214 101754 4220 101756
rect 4276 101754 4300 101756
rect 4356 101754 4380 101756
rect 4436 101754 4460 101756
rect 4516 101754 4522 101756
rect 4276 101702 4278 101754
rect 4458 101702 4460 101754
rect 4214 101700 4220 101702
rect 4276 101700 4300 101702
rect 4356 101700 4380 101702
rect 4436 101700 4460 101702
rect 4516 101700 4522 101702
rect 4214 101680 4522 101700
rect 4214 100668 4522 100688
rect 4214 100666 4220 100668
rect 4276 100666 4300 100668
rect 4356 100666 4380 100668
rect 4436 100666 4460 100668
rect 4516 100666 4522 100668
rect 4276 100614 4278 100666
rect 4458 100614 4460 100666
rect 4214 100612 4220 100614
rect 4276 100612 4300 100614
rect 4356 100612 4380 100614
rect 4436 100612 4460 100614
rect 4516 100612 4522 100614
rect 4214 100592 4522 100612
rect 4214 99580 4522 99600
rect 4214 99578 4220 99580
rect 4276 99578 4300 99580
rect 4356 99578 4380 99580
rect 4436 99578 4460 99580
rect 4516 99578 4522 99580
rect 4276 99526 4278 99578
rect 4458 99526 4460 99578
rect 4214 99524 4220 99526
rect 4276 99524 4300 99526
rect 4356 99524 4380 99526
rect 4436 99524 4460 99526
rect 4516 99524 4522 99526
rect 4214 99504 4522 99524
rect 4214 98492 4522 98512
rect 4214 98490 4220 98492
rect 4276 98490 4300 98492
rect 4356 98490 4380 98492
rect 4436 98490 4460 98492
rect 4516 98490 4522 98492
rect 4276 98438 4278 98490
rect 4458 98438 4460 98490
rect 4214 98436 4220 98438
rect 4276 98436 4300 98438
rect 4356 98436 4380 98438
rect 4436 98436 4460 98438
rect 4516 98436 4522 98438
rect 4214 98416 4522 98436
rect 4214 97404 4522 97424
rect 4214 97402 4220 97404
rect 4276 97402 4300 97404
rect 4356 97402 4380 97404
rect 4436 97402 4460 97404
rect 4516 97402 4522 97404
rect 4276 97350 4278 97402
rect 4458 97350 4460 97402
rect 4214 97348 4220 97350
rect 4276 97348 4300 97350
rect 4356 97348 4380 97350
rect 4436 97348 4460 97350
rect 4516 97348 4522 97350
rect 4214 97328 4522 97348
rect 4214 96316 4522 96336
rect 4214 96314 4220 96316
rect 4276 96314 4300 96316
rect 4356 96314 4380 96316
rect 4436 96314 4460 96316
rect 4516 96314 4522 96316
rect 4276 96262 4278 96314
rect 4458 96262 4460 96314
rect 4214 96260 4220 96262
rect 4276 96260 4300 96262
rect 4356 96260 4380 96262
rect 4436 96260 4460 96262
rect 4516 96260 4522 96262
rect 4214 96240 4522 96260
rect 4214 95228 4522 95248
rect 4214 95226 4220 95228
rect 4276 95226 4300 95228
rect 4356 95226 4380 95228
rect 4436 95226 4460 95228
rect 4516 95226 4522 95228
rect 4276 95174 4278 95226
rect 4458 95174 4460 95226
rect 4214 95172 4220 95174
rect 4276 95172 4300 95174
rect 4356 95172 4380 95174
rect 4436 95172 4460 95174
rect 4516 95172 4522 95174
rect 4214 95152 4522 95172
rect 2964 94444 3016 94450
rect 2964 94386 3016 94392
rect 2780 79212 2832 79218
rect 2780 79154 2832 79160
rect 2596 78600 2648 78606
rect 2596 78542 2648 78548
rect 2608 78266 2636 78542
rect 2596 78260 2648 78266
rect 2596 78202 2648 78208
rect 2792 78130 2820 79154
rect 2780 78124 2832 78130
rect 2780 78066 2832 78072
rect 2320 66156 2372 66162
rect 2320 66098 2372 66104
rect 2332 65550 2360 66098
rect 2320 65544 2372 65550
rect 2320 65486 2372 65492
rect 2228 60104 2280 60110
rect 2228 60046 2280 60052
rect 1952 59628 2004 59634
rect 1952 59570 2004 59576
rect 2976 59226 3004 94386
rect 4214 94140 4522 94160
rect 4214 94138 4220 94140
rect 4276 94138 4300 94140
rect 4356 94138 4380 94140
rect 4436 94138 4460 94140
rect 4516 94138 4522 94140
rect 4276 94086 4278 94138
rect 4458 94086 4460 94138
rect 4214 94084 4220 94086
rect 4276 94084 4300 94086
rect 4356 94084 4380 94086
rect 4436 94084 4460 94086
rect 4516 94084 4522 94086
rect 4214 94064 4522 94084
rect 4214 93052 4522 93072
rect 4214 93050 4220 93052
rect 4276 93050 4300 93052
rect 4356 93050 4380 93052
rect 4436 93050 4460 93052
rect 4516 93050 4522 93052
rect 4276 92998 4278 93050
rect 4458 92998 4460 93050
rect 4214 92996 4220 92998
rect 4276 92996 4300 92998
rect 4356 92996 4380 92998
rect 4436 92996 4460 92998
rect 4516 92996 4522 92998
rect 4214 92976 4522 92996
rect 4214 91964 4522 91984
rect 4214 91962 4220 91964
rect 4276 91962 4300 91964
rect 4356 91962 4380 91964
rect 4436 91962 4460 91964
rect 4516 91962 4522 91964
rect 4276 91910 4278 91962
rect 4458 91910 4460 91962
rect 4214 91908 4220 91910
rect 4276 91908 4300 91910
rect 4356 91908 4380 91910
rect 4436 91908 4460 91910
rect 4516 91908 4522 91910
rect 4214 91888 4522 91908
rect 4214 90876 4522 90896
rect 4214 90874 4220 90876
rect 4276 90874 4300 90876
rect 4356 90874 4380 90876
rect 4436 90874 4460 90876
rect 4516 90874 4522 90876
rect 4276 90822 4278 90874
rect 4458 90822 4460 90874
rect 4214 90820 4220 90822
rect 4276 90820 4300 90822
rect 4356 90820 4380 90822
rect 4436 90820 4460 90822
rect 4516 90820 4522 90822
rect 4214 90800 4522 90820
rect 4214 89788 4522 89808
rect 4214 89786 4220 89788
rect 4276 89786 4300 89788
rect 4356 89786 4380 89788
rect 4436 89786 4460 89788
rect 4516 89786 4522 89788
rect 4276 89734 4278 89786
rect 4458 89734 4460 89786
rect 4214 89732 4220 89734
rect 4276 89732 4300 89734
rect 4356 89732 4380 89734
rect 4436 89732 4460 89734
rect 4516 89732 4522 89734
rect 4214 89712 4522 89732
rect 7852 88806 7880 117234
rect 8036 117094 8064 119326
rect 11610 119326 11744 119354
rect 11610 119200 11666 119326
rect 11716 117298 11744 119326
rect 15474 119326 15792 119354
rect 15474 119200 15530 119326
rect 11704 117292 11756 117298
rect 11704 117234 11756 117240
rect 15568 117292 15620 117298
rect 15568 117234 15620 117240
rect 11888 117224 11940 117230
rect 11888 117166 11940 117172
rect 8024 117088 8076 117094
rect 8024 117030 8076 117036
rect 10692 116816 10744 116822
rect 10692 116758 10744 116764
rect 7840 88800 7892 88806
rect 7840 88742 7892 88748
rect 4214 88700 4522 88720
rect 4214 88698 4220 88700
rect 4276 88698 4300 88700
rect 4356 88698 4380 88700
rect 4436 88698 4460 88700
rect 4516 88698 4522 88700
rect 4276 88646 4278 88698
rect 4458 88646 4460 88698
rect 4214 88644 4220 88646
rect 4276 88644 4300 88646
rect 4356 88644 4380 88646
rect 4436 88644 4460 88646
rect 4516 88644 4522 88646
rect 4214 88624 4522 88644
rect 4214 87612 4522 87632
rect 4214 87610 4220 87612
rect 4276 87610 4300 87612
rect 4356 87610 4380 87612
rect 4436 87610 4460 87612
rect 4516 87610 4522 87612
rect 4276 87558 4278 87610
rect 4458 87558 4460 87610
rect 4214 87556 4220 87558
rect 4276 87556 4300 87558
rect 4356 87556 4380 87558
rect 4436 87556 4460 87558
rect 4516 87556 4522 87558
rect 4214 87536 4522 87556
rect 4214 86524 4522 86544
rect 4214 86522 4220 86524
rect 4276 86522 4300 86524
rect 4356 86522 4380 86524
rect 4436 86522 4460 86524
rect 4516 86522 4522 86524
rect 4276 86470 4278 86522
rect 4458 86470 4460 86522
rect 4214 86468 4220 86470
rect 4276 86468 4300 86470
rect 4356 86468 4380 86470
rect 4436 86468 4460 86470
rect 4516 86468 4522 86470
rect 4214 86448 4522 86468
rect 4214 85436 4522 85456
rect 4214 85434 4220 85436
rect 4276 85434 4300 85436
rect 4356 85434 4380 85436
rect 4436 85434 4460 85436
rect 4516 85434 4522 85436
rect 4276 85382 4278 85434
rect 4458 85382 4460 85434
rect 4214 85380 4220 85382
rect 4276 85380 4300 85382
rect 4356 85380 4380 85382
rect 4436 85380 4460 85382
rect 4516 85380 4522 85382
rect 4214 85360 4522 85380
rect 4214 84348 4522 84368
rect 4214 84346 4220 84348
rect 4276 84346 4300 84348
rect 4356 84346 4380 84348
rect 4436 84346 4460 84348
rect 4516 84346 4522 84348
rect 4276 84294 4278 84346
rect 4458 84294 4460 84346
rect 4214 84292 4220 84294
rect 4276 84292 4300 84294
rect 4356 84292 4380 84294
rect 4436 84292 4460 84294
rect 4516 84292 4522 84294
rect 4214 84272 4522 84292
rect 4214 83260 4522 83280
rect 4214 83258 4220 83260
rect 4276 83258 4300 83260
rect 4356 83258 4380 83260
rect 4436 83258 4460 83260
rect 4516 83258 4522 83260
rect 4276 83206 4278 83258
rect 4458 83206 4460 83258
rect 4214 83204 4220 83206
rect 4276 83204 4300 83206
rect 4356 83204 4380 83206
rect 4436 83204 4460 83206
rect 4516 83204 4522 83206
rect 4214 83184 4522 83204
rect 4214 82172 4522 82192
rect 4214 82170 4220 82172
rect 4276 82170 4300 82172
rect 4356 82170 4380 82172
rect 4436 82170 4460 82172
rect 4516 82170 4522 82172
rect 4276 82118 4278 82170
rect 4458 82118 4460 82170
rect 4214 82116 4220 82118
rect 4276 82116 4300 82118
rect 4356 82116 4380 82118
rect 4436 82116 4460 82118
rect 4516 82116 4522 82118
rect 4214 82096 4522 82116
rect 4214 81084 4522 81104
rect 4214 81082 4220 81084
rect 4276 81082 4300 81084
rect 4356 81082 4380 81084
rect 4436 81082 4460 81084
rect 4516 81082 4522 81084
rect 4276 81030 4278 81082
rect 4458 81030 4460 81082
rect 4214 81028 4220 81030
rect 4276 81028 4300 81030
rect 4356 81028 4380 81030
rect 4436 81028 4460 81030
rect 4516 81028 4522 81030
rect 4214 81008 4522 81028
rect 4214 79996 4522 80016
rect 4214 79994 4220 79996
rect 4276 79994 4300 79996
rect 4356 79994 4380 79996
rect 4436 79994 4460 79996
rect 4516 79994 4522 79996
rect 4276 79942 4278 79994
rect 4458 79942 4460 79994
rect 4214 79940 4220 79942
rect 4276 79940 4300 79942
rect 4356 79940 4380 79942
rect 4436 79940 4460 79942
rect 4516 79940 4522 79942
rect 4214 79920 4522 79940
rect 10704 79354 10732 116758
rect 10692 79348 10744 79354
rect 10692 79290 10744 79296
rect 4214 78908 4522 78928
rect 4214 78906 4220 78908
rect 4276 78906 4300 78908
rect 4356 78906 4380 78908
rect 4436 78906 4460 78908
rect 4516 78906 4522 78908
rect 4276 78854 4278 78906
rect 4458 78854 4460 78906
rect 4214 78852 4220 78854
rect 4276 78852 4300 78854
rect 4356 78852 4380 78854
rect 4436 78852 4460 78854
rect 4516 78852 4522 78854
rect 4214 78832 4522 78852
rect 3056 78124 3108 78130
rect 3056 78066 3108 78072
rect 2964 59220 3016 59226
rect 2964 59162 3016 59168
rect 2964 59016 3016 59022
rect 2964 58958 3016 58964
rect 2976 58546 3004 58958
rect 2964 58540 3016 58546
rect 2964 58482 3016 58488
rect 1412 55186 1532 55214
rect 1596 58398 1808 58426
rect 1412 31906 1440 55186
rect 1492 54528 1544 54534
rect 1490 54496 1492 54505
rect 1544 54496 1546 54505
rect 1490 54431 1546 54440
rect 1492 50720 1544 50726
rect 1492 50662 1544 50668
rect 1504 50425 1532 50662
rect 1490 50416 1546 50425
rect 1490 50351 1546 50360
rect 1596 50266 1624 58398
rect 1676 58336 1728 58342
rect 1676 58278 1728 58284
rect 1504 50238 1624 50266
rect 1504 35086 1532 50238
rect 1584 47184 1636 47190
rect 1584 47126 1636 47132
rect 1596 47025 1624 47126
rect 1582 47016 1638 47025
rect 1582 46951 1638 46960
rect 1492 35080 1544 35086
rect 1492 35022 1544 35028
rect 1584 34944 1636 34950
rect 1584 34886 1636 34892
rect 1596 34785 1624 34886
rect 1582 34776 1638 34785
rect 1582 34711 1638 34720
rect 1412 31878 1532 31906
rect 1400 31816 1452 31822
rect 1400 31758 1452 31764
rect 1412 31385 1440 31758
rect 1398 31376 1454 31385
rect 1398 31311 1454 31320
rect 1400 27464 1452 27470
rect 1400 27406 1452 27412
rect 1412 27305 1440 27406
rect 1398 27296 1454 27305
rect 1398 27231 1454 27240
rect 1400 23724 1452 23730
rect 1400 23666 1452 23672
rect 1412 23225 1440 23666
rect 1398 23216 1454 23225
rect 1398 23151 1454 23160
rect 1504 19378 1532 31878
rect 1492 19372 1544 19378
rect 1492 19314 1544 19320
rect 1584 19168 1636 19174
rect 1582 19136 1584 19145
rect 1636 19136 1638 19145
rect 1582 19071 1638 19080
rect 1492 15904 1544 15910
rect 1492 15846 1544 15852
rect 1504 15745 1532 15846
rect 1490 15736 1546 15745
rect 1490 15671 1546 15680
rect 1400 11756 1452 11762
rect 1400 11698 1452 11704
rect 1412 11665 1440 11698
rect 1398 11656 1454 11665
rect 1398 11591 1454 11600
rect 1584 7744 1636 7750
rect 1584 7686 1636 7692
rect 1596 7585 1624 7686
rect 1582 7576 1638 7585
rect 1582 7511 1638 7520
rect 1688 3602 1716 58278
rect 2872 47048 2924 47054
rect 2872 46990 2924 46996
rect 1860 43308 1912 43314
rect 1860 43250 1912 43256
rect 1872 42945 1900 43250
rect 1858 42936 1914 42945
rect 1858 42871 1914 42880
rect 1860 38956 1912 38962
rect 1860 38898 1912 38904
rect 1872 38865 1900 38898
rect 1858 38856 1914 38865
rect 1858 38791 1914 38800
rect 1768 25492 1820 25498
rect 1768 25434 1820 25440
rect 1780 16250 1808 25434
rect 1768 16244 1820 16250
rect 1768 16186 1820 16192
rect 2884 13530 2912 46990
rect 2872 13524 2924 13530
rect 2872 13466 2924 13472
rect 2412 13320 2464 13326
rect 2412 13262 2464 13268
rect 2424 7546 2452 13262
rect 2688 7880 2740 7886
rect 2688 7822 2740 7828
rect 2700 7546 2728 7822
rect 2412 7540 2464 7546
rect 2412 7482 2464 7488
rect 2688 7540 2740 7546
rect 2688 7482 2740 7488
rect 1676 3596 1728 3602
rect 1676 3538 1728 3544
rect 1400 3528 1452 3534
rect 1398 3496 1400 3505
rect 1452 3496 1454 3505
rect 1398 3431 1454 3440
rect 20 2440 72 2446
rect 20 2382 72 2388
rect 32 800 60 2382
rect 2976 2038 3004 58482
rect 3068 11830 3096 78066
rect 4214 77820 4522 77840
rect 4214 77818 4220 77820
rect 4276 77818 4300 77820
rect 4356 77818 4380 77820
rect 4436 77818 4460 77820
rect 4516 77818 4522 77820
rect 4276 77766 4278 77818
rect 4458 77766 4460 77818
rect 4214 77764 4220 77766
rect 4276 77764 4300 77766
rect 4356 77764 4380 77766
rect 4436 77764 4460 77766
rect 4516 77764 4522 77766
rect 4214 77744 4522 77764
rect 4214 76732 4522 76752
rect 4214 76730 4220 76732
rect 4276 76730 4300 76732
rect 4356 76730 4380 76732
rect 4436 76730 4460 76732
rect 4516 76730 4522 76732
rect 4276 76678 4278 76730
rect 4458 76678 4460 76730
rect 4214 76676 4220 76678
rect 4276 76676 4300 76678
rect 4356 76676 4380 76678
rect 4436 76676 4460 76678
rect 4516 76676 4522 76678
rect 4214 76656 4522 76676
rect 4214 75644 4522 75664
rect 4214 75642 4220 75644
rect 4276 75642 4300 75644
rect 4356 75642 4380 75644
rect 4436 75642 4460 75644
rect 4516 75642 4522 75644
rect 4276 75590 4278 75642
rect 4458 75590 4460 75642
rect 4214 75588 4220 75590
rect 4276 75588 4300 75590
rect 4356 75588 4380 75590
rect 4436 75588 4460 75590
rect 4516 75588 4522 75590
rect 4214 75568 4522 75588
rect 4214 74556 4522 74576
rect 4214 74554 4220 74556
rect 4276 74554 4300 74556
rect 4356 74554 4380 74556
rect 4436 74554 4460 74556
rect 4516 74554 4522 74556
rect 4276 74502 4278 74554
rect 4458 74502 4460 74554
rect 4214 74500 4220 74502
rect 4276 74500 4300 74502
rect 4356 74500 4380 74502
rect 4436 74500 4460 74502
rect 4516 74500 4522 74502
rect 4214 74480 4522 74500
rect 4214 73468 4522 73488
rect 4214 73466 4220 73468
rect 4276 73466 4300 73468
rect 4356 73466 4380 73468
rect 4436 73466 4460 73468
rect 4516 73466 4522 73468
rect 4276 73414 4278 73466
rect 4458 73414 4460 73466
rect 4214 73412 4220 73414
rect 4276 73412 4300 73414
rect 4356 73412 4380 73414
rect 4436 73412 4460 73414
rect 4516 73412 4522 73414
rect 4214 73392 4522 73412
rect 4214 72380 4522 72400
rect 4214 72378 4220 72380
rect 4276 72378 4300 72380
rect 4356 72378 4380 72380
rect 4436 72378 4460 72380
rect 4516 72378 4522 72380
rect 4276 72326 4278 72378
rect 4458 72326 4460 72378
rect 4214 72324 4220 72326
rect 4276 72324 4300 72326
rect 4356 72324 4380 72326
rect 4436 72324 4460 72326
rect 4516 72324 4522 72326
rect 4214 72304 4522 72324
rect 4214 71292 4522 71312
rect 4214 71290 4220 71292
rect 4276 71290 4300 71292
rect 4356 71290 4380 71292
rect 4436 71290 4460 71292
rect 4516 71290 4522 71292
rect 4276 71238 4278 71290
rect 4458 71238 4460 71290
rect 4214 71236 4220 71238
rect 4276 71236 4300 71238
rect 4356 71236 4380 71238
rect 4436 71236 4460 71238
rect 4516 71236 4522 71238
rect 4214 71216 4522 71236
rect 4214 70204 4522 70224
rect 4214 70202 4220 70204
rect 4276 70202 4300 70204
rect 4356 70202 4380 70204
rect 4436 70202 4460 70204
rect 4516 70202 4522 70204
rect 4276 70150 4278 70202
rect 4458 70150 4460 70202
rect 4214 70148 4220 70150
rect 4276 70148 4300 70150
rect 4356 70148 4380 70150
rect 4436 70148 4460 70150
rect 4516 70148 4522 70150
rect 4214 70128 4522 70148
rect 4214 69116 4522 69136
rect 4214 69114 4220 69116
rect 4276 69114 4300 69116
rect 4356 69114 4380 69116
rect 4436 69114 4460 69116
rect 4516 69114 4522 69116
rect 4276 69062 4278 69114
rect 4458 69062 4460 69114
rect 4214 69060 4220 69062
rect 4276 69060 4300 69062
rect 4356 69060 4380 69062
rect 4436 69060 4460 69062
rect 4516 69060 4522 69062
rect 4214 69040 4522 69060
rect 4214 68028 4522 68048
rect 4214 68026 4220 68028
rect 4276 68026 4300 68028
rect 4356 68026 4380 68028
rect 4436 68026 4460 68028
rect 4516 68026 4522 68028
rect 4276 67974 4278 68026
rect 4458 67974 4460 68026
rect 4214 67972 4220 67974
rect 4276 67972 4300 67974
rect 4356 67972 4380 67974
rect 4436 67972 4460 67974
rect 4516 67972 4522 67974
rect 4214 67952 4522 67972
rect 4214 66940 4522 66960
rect 4214 66938 4220 66940
rect 4276 66938 4300 66940
rect 4356 66938 4380 66940
rect 4436 66938 4460 66940
rect 4516 66938 4522 66940
rect 4276 66886 4278 66938
rect 4458 66886 4460 66938
rect 4214 66884 4220 66886
rect 4276 66884 4300 66886
rect 4356 66884 4380 66886
rect 4436 66884 4460 66886
rect 4516 66884 4522 66886
rect 4214 66864 4522 66884
rect 4214 65852 4522 65872
rect 4214 65850 4220 65852
rect 4276 65850 4300 65852
rect 4356 65850 4380 65852
rect 4436 65850 4460 65852
rect 4516 65850 4522 65852
rect 4276 65798 4278 65850
rect 4458 65798 4460 65850
rect 4214 65796 4220 65798
rect 4276 65796 4300 65798
rect 4356 65796 4380 65798
rect 4436 65796 4460 65798
rect 4516 65796 4522 65798
rect 4214 65776 4522 65796
rect 11900 65482 11928 117166
rect 15580 116890 15608 117234
rect 15764 117094 15792 119326
rect 19338 119200 19394 120000
rect 22558 119354 22614 120000
rect 22558 119326 22876 119354
rect 22558 119200 22614 119326
rect 19352 117162 19380 119200
rect 19574 117532 19882 117552
rect 19574 117530 19580 117532
rect 19636 117530 19660 117532
rect 19716 117530 19740 117532
rect 19796 117530 19820 117532
rect 19876 117530 19882 117532
rect 19636 117478 19638 117530
rect 19818 117478 19820 117530
rect 19574 117476 19580 117478
rect 19636 117476 19660 117478
rect 19716 117476 19740 117478
rect 19796 117476 19820 117478
rect 19876 117476 19882 117478
rect 19574 117456 19882 117476
rect 19432 117292 19484 117298
rect 19432 117234 19484 117240
rect 22652 117292 22704 117298
rect 22652 117234 22704 117240
rect 19340 117156 19392 117162
rect 19340 117098 19392 117104
rect 15752 117088 15804 117094
rect 15752 117030 15804 117036
rect 15568 116884 15620 116890
rect 15568 116826 15620 116832
rect 11888 65476 11940 65482
rect 11888 65418 11940 65424
rect 4214 64764 4522 64784
rect 4214 64762 4220 64764
rect 4276 64762 4300 64764
rect 4356 64762 4380 64764
rect 4436 64762 4460 64764
rect 4516 64762 4522 64764
rect 4276 64710 4278 64762
rect 4458 64710 4460 64762
rect 4214 64708 4220 64710
rect 4276 64708 4300 64710
rect 4356 64708 4380 64710
rect 4436 64708 4460 64710
rect 4516 64708 4522 64710
rect 4214 64688 4522 64708
rect 4214 63676 4522 63696
rect 4214 63674 4220 63676
rect 4276 63674 4300 63676
rect 4356 63674 4380 63676
rect 4436 63674 4460 63676
rect 4516 63674 4522 63676
rect 4276 63622 4278 63674
rect 4458 63622 4460 63674
rect 4214 63620 4220 63622
rect 4276 63620 4300 63622
rect 4356 63620 4380 63622
rect 4436 63620 4460 63622
rect 4516 63620 4522 63622
rect 4214 63600 4522 63620
rect 4214 62588 4522 62608
rect 4214 62586 4220 62588
rect 4276 62586 4300 62588
rect 4356 62586 4380 62588
rect 4436 62586 4460 62588
rect 4516 62586 4522 62588
rect 4276 62534 4278 62586
rect 4458 62534 4460 62586
rect 4214 62532 4220 62534
rect 4276 62532 4300 62534
rect 4356 62532 4380 62534
rect 4436 62532 4460 62534
rect 4516 62532 4522 62534
rect 4214 62512 4522 62532
rect 4214 61500 4522 61520
rect 4214 61498 4220 61500
rect 4276 61498 4300 61500
rect 4356 61498 4380 61500
rect 4436 61498 4460 61500
rect 4516 61498 4522 61500
rect 4276 61446 4278 61498
rect 4458 61446 4460 61498
rect 4214 61444 4220 61446
rect 4276 61444 4300 61446
rect 4356 61444 4380 61446
rect 4436 61444 4460 61446
rect 4516 61444 4522 61446
rect 4214 61424 4522 61444
rect 19444 61130 19472 117234
rect 19574 116444 19882 116464
rect 19574 116442 19580 116444
rect 19636 116442 19660 116444
rect 19716 116442 19740 116444
rect 19796 116442 19820 116444
rect 19876 116442 19882 116444
rect 19636 116390 19638 116442
rect 19818 116390 19820 116442
rect 19574 116388 19580 116390
rect 19636 116388 19660 116390
rect 19716 116388 19740 116390
rect 19796 116388 19820 116390
rect 19876 116388 19882 116390
rect 19574 116368 19882 116388
rect 19574 115356 19882 115376
rect 19574 115354 19580 115356
rect 19636 115354 19660 115356
rect 19716 115354 19740 115356
rect 19796 115354 19820 115356
rect 19876 115354 19882 115356
rect 19636 115302 19638 115354
rect 19818 115302 19820 115354
rect 19574 115300 19580 115302
rect 19636 115300 19660 115302
rect 19716 115300 19740 115302
rect 19796 115300 19820 115302
rect 19876 115300 19882 115302
rect 19574 115280 19882 115300
rect 19574 114268 19882 114288
rect 19574 114266 19580 114268
rect 19636 114266 19660 114268
rect 19716 114266 19740 114268
rect 19796 114266 19820 114268
rect 19876 114266 19882 114268
rect 19636 114214 19638 114266
rect 19818 114214 19820 114266
rect 19574 114212 19580 114214
rect 19636 114212 19660 114214
rect 19716 114212 19740 114214
rect 19796 114212 19820 114214
rect 19876 114212 19882 114214
rect 19574 114192 19882 114212
rect 20628 114028 20680 114034
rect 20628 113970 20680 113976
rect 19574 113180 19882 113200
rect 19574 113178 19580 113180
rect 19636 113178 19660 113180
rect 19716 113178 19740 113180
rect 19796 113178 19820 113180
rect 19876 113178 19882 113180
rect 19636 113126 19638 113178
rect 19818 113126 19820 113178
rect 19574 113124 19580 113126
rect 19636 113124 19660 113126
rect 19716 113124 19740 113126
rect 19796 113124 19820 113126
rect 19876 113124 19882 113126
rect 19574 113104 19882 113124
rect 19574 112092 19882 112112
rect 19574 112090 19580 112092
rect 19636 112090 19660 112092
rect 19716 112090 19740 112092
rect 19796 112090 19820 112092
rect 19876 112090 19882 112092
rect 19636 112038 19638 112090
rect 19818 112038 19820 112090
rect 19574 112036 19580 112038
rect 19636 112036 19660 112038
rect 19716 112036 19740 112038
rect 19796 112036 19820 112038
rect 19876 112036 19882 112038
rect 19574 112016 19882 112036
rect 19574 111004 19882 111024
rect 19574 111002 19580 111004
rect 19636 111002 19660 111004
rect 19716 111002 19740 111004
rect 19796 111002 19820 111004
rect 19876 111002 19882 111004
rect 19636 110950 19638 111002
rect 19818 110950 19820 111002
rect 19574 110948 19580 110950
rect 19636 110948 19660 110950
rect 19716 110948 19740 110950
rect 19796 110948 19820 110950
rect 19876 110948 19882 110950
rect 19574 110928 19882 110948
rect 19574 109916 19882 109936
rect 19574 109914 19580 109916
rect 19636 109914 19660 109916
rect 19716 109914 19740 109916
rect 19796 109914 19820 109916
rect 19876 109914 19882 109916
rect 19636 109862 19638 109914
rect 19818 109862 19820 109914
rect 19574 109860 19580 109862
rect 19636 109860 19660 109862
rect 19716 109860 19740 109862
rect 19796 109860 19820 109862
rect 19876 109860 19882 109862
rect 19574 109840 19882 109860
rect 20640 109478 20668 113970
rect 20628 109472 20680 109478
rect 20628 109414 20680 109420
rect 19574 108828 19882 108848
rect 19574 108826 19580 108828
rect 19636 108826 19660 108828
rect 19716 108826 19740 108828
rect 19796 108826 19820 108828
rect 19876 108826 19882 108828
rect 19636 108774 19638 108826
rect 19818 108774 19820 108826
rect 19574 108772 19580 108774
rect 19636 108772 19660 108774
rect 19716 108772 19740 108774
rect 19796 108772 19820 108774
rect 19876 108772 19882 108774
rect 19574 108752 19882 108772
rect 19574 107740 19882 107760
rect 19574 107738 19580 107740
rect 19636 107738 19660 107740
rect 19716 107738 19740 107740
rect 19796 107738 19820 107740
rect 19876 107738 19882 107740
rect 19636 107686 19638 107738
rect 19818 107686 19820 107738
rect 19574 107684 19580 107686
rect 19636 107684 19660 107686
rect 19716 107684 19740 107686
rect 19796 107684 19820 107686
rect 19876 107684 19882 107686
rect 19574 107664 19882 107684
rect 19574 106652 19882 106672
rect 19574 106650 19580 106652
rect 19636 106650 19660 106652
rect 19716 106650 19740 106652
rect 19796 106650 19820 106652
rect 19876 106650 19882 106652
rect 19636 106598 19638 106650
rect 19818 106598 19820 106650
rect 19574 106596 19580 106598
rect 19636 106596 19660 106598
rect 19716 106596 19740 106598
rect 19796 106596 19820 106598
rect 19876 106596 19882 106598
rect 19574 106576 19882 106596
rect 19574 105564 19882 105584
rect 19574 105562 19580 105564
rect 19636 105562 19660 105564
rect 19716 105562 19740 105564
rect 19796 105562 19820 105564
rect 19876 105562 19882 105564
rect 19636 105510 19638 105562
rect 19818 105510 19820 105562
rect 19574 105508 19580 105510
rect 19636 105508 19660 105510
rect 19716 105508 19740 105510
rect 19796 105508 19820 105510
rect 19876 105508 19882 105510
rect 19574 105488 19882 105508
rect 19574 104476 19882 104496
rect 19574 104474 19580 104476
rect 19636 104474 19660 104476
rect 19716 104474 19740 104476
rect 19796 104474 19820 104476
rect 19876 104474 19882 104476
rect 19636 104422 19638 104474
rect 19818 104422 19820 104474
rect 19574 104420 19580 104422
rect 19636 104420 19660 104422
rect 19716 104420 19740 104422
rect 19796 104420 19820 104422
rect 19876 104420 19882 104422
rect 19574 104400 19882 104420
rect 19574 103388 19882 103408
rect 19574 103386 19580 103388
rect 19636 103386 19660 103388
rect 19716 103386 19740 103388
rect 19796 103386 19820 103388
rect 19876 103386 19882 103388
rect 19636 103334 19638 103386
rect 19818 103334 19820 103386
rect 19574 103332 19580 103334
rect 19636 103332 19660 103334
rect 19716 103332 19740 103334
rect 19796 103332 19820 103334
rect 19876 103332 19882 103334
rect 19574 103312 19882 103332
rect 19574 102300 19882 102320
rect 19574 102298 19580 102300
rect 19636 102298 19660 102300
rect 19716 102298 19740 102300
rect 19796 102298 19820 102300
rect 19876 102298 19882 102300
rect 19636 102246 19638 102298
rect 19818 102246 19820 102298
rect 19574 102244 19580 102246
rect 19636 102244 19660 102246
rect 19716 102244 19740 102246
rect 19796 102244 19820 102246
rect 19876 102244 19882 102246
rect 19574 102224 19882 102244
rect 19574 101212 19882 101232
rect 19574 101210 19580 101212
rect 19636 101210 19660 101212
rect 19716 101210 19740 101212
rect 19796 101210 19820 101212
rect 19876 101210 19882 101212
rect 19636 101158 19638 101210
rect 19818 101158 19820 101210
rect 19574 101156 19580 101158
rect 19636 101156 19660 101158
rect 19716 101156 19740 101158
rect 19796 101156 19820 101158
rect 19876 101156 19882 101158
rect 19574 101136 19882 101156
rect 19574 100124 19882 100144
rect 19574 100122 19580 100124
rect 19636 100122 19660 100124
rect 19716 100122 19740 100124
rect 19796 100122 19820 100124
rect 19876 100122 19882 100124
rect 19636 100070 19638 100122
rect 19818 100070 19820 100122
rect 19574 100068 19580 100070
rect 19636 100068 19660 100070
rect 19716 100068 19740 100070
rect 19796 100068 19820 100070
rect 19876 100068 19882 100070
rect 19574 100048 19882 100068
rect 19574 99036 19882 99056
rect 19574 99034 19580 99036
rect 19636 99034 19660 99036
rect 19716 99034 19740 99036
rect 19796 99034 19820 99036
rect 19876 99034 19882 99036
rect 19636 98982 19638 99034
rect 19818 98982 19820 99034
rect 19574 98980 19580 98982
rect 19636 98980 19660 98982
rect 19716 98980 19740 98982
rect 19796 98980 19820 98982
rect 19876 98980 19882 98982
rect 19574 98960 19882 98980
rect 19574 97948 19882 97968
rect 19574 97946 19580 97948
rect 19636 97946 19660 97948
rect 19716 97946 19740 97948
rect 19796 97946 19820 97948
rect 19876 97946 19882 97948
rect 19636 97894 19638 97946
rect 19818 97894 19820 97946
rect 19574 97892 19580 97894
rect 19636 97892 19660 97894
rect 19716 97892 19740 97894
rect 19796 97892 19820 97894
rect 19876 97892 19882 97894
rect 19574 97872 19882 97892
rect 19574 96860 19882 96880
rect 19574 96858 19580 96860
rect 19636 96858 19660 96860
rect 19716 96858 19740 96860
rect 19796 96858 19820 96860
rect 19876 96858 19882 96860
rect 19636 96806 19638 96858
rect 19818 96806 19820 96858
rect 19574 96804 19580 96806
rect 19636 96804 19660 96806
rect 19716 96804 19740 96806
rect 19796 96804 19820 96806
rect 19876 96804 19882 96806
rect 19574 96784 19882 96804
rect 19574 95772 19882 95792
rect 19574 95770 19580 95772
rect 19636 95770 19660 95772
rect 19716 95770 19740 95772
rect 19796 95770 19820 95772
rect 19876 95770 19882 95772
rect 19636 95718 19638 95770
rect 19818 95718 19820 95770
rect 19574 95716 19580 95718
rect 19636 95716 19660 95718
rect 19716 95716 19740 95718
rect 19796 95716 19820 95718
rect 19876 95716 19882 95718
rect 19574 95696 19882 95716
rect 19574 94684 19882 94704
rect 19574 94682 19580 94684
rect 19636 94682 19660 94684
rect 19716 94682 19740 94684
rect 19796 94682 19820 94684
rect 19876 94682 19882 94684
rect 19636 94630 19638 94682
rect 19818 94630 19820 94682
rect 19574 94628 19580 94630
rect 19636 94628 19660 94630
rect 19716 94628 19740 94630
rect 19796 94628 19820 94630
rect 19876 94628 19882 94630
rect 19574 94608 19882 94628
rect 19574 93596 19882 93616
rect 19574 93594 19580 93596
rect 19636 93594 19660 93596
rect 19716 93594 19740 93596
rect 19796 93594 19820 93596
rect 19876 93594 19882 93596
rect 19636 93542 19638 93594
rect 19818 93542 19820 93594
rect 19574 93540 19580 93542
rect 19636 93540 19660 93542
rect 19716 93540 19740 93542
rect 19796 93540 19820 93542
rect 19876 93540 19882 93542
rect 19574 93520 19882 93540
rect 19574 92508 19882 92528
rect 19574 92506 19580 92508
rect 19636 92506 19660 92508
rect 19716 92506 19740 92508
rect 19796 92506 19820 92508
rect 19876 92506 19882 92508
rect 19636 92454 19638 92506
rect 19818 92454 19820 92506
rect 19574 92452 19580 92454
rect 19636 92452 19660 92454
rect 19716 92452 19740 92454
rect 19796 92452 19820 92454
rect 19876 92452 19882 92454
rect 19574 92432 19882 92452
rect 19574 91420 19882 91440
rect 19574 91418 19580 91420
rect 19636 91418 19660 91420
rect 19716 91418 19740 91420
rect 19796 91418 19820 91420
rect 19876 91418 19882 91420
rect 19636 91366 19638 91418
rect 19818 91366 19820 91418
rect 19574 91364 19580 91366
rect 19636 91364 19660 91366
rect 19716 91364 19740 91366
rect 19796 91364 19820 91366
rect 19876 91364 19882 91366
rect 19574 91344 19882 91364
rect 19574 90332 19882 90352
rect 19574 90330 19580 90332
rect 19636 90330 19660 90332
rect 19716 90330 19740 90332
rect 19796 90330 19820 90332
rect 19876 90330 19882 90332
rect 19636 90278 19638 90330
rect 19818 90278 19820 90330
rect 19574 90276 19580 90278
rect 19636 90276 19660 90278
rect 19716 90276 19740 90278
rect 19796 90276 19820 90278
rect 19876 90276 19882 90278
rect 19574 90256 19882 90276
rect 19574 89244 19882 89264
rect 19574 89242 19580 89244
rect 19636 89242 19660 89244
rect 19716 89242 19740 89244
rect 19796 89242 19820 89244
rect 19876 89242 19882 89244
rect 19636 89190 19638 89242
rect 19818 89190 19820 89242
rect 19574 89188 19580 89190
rect 19636 89188 19660 89190
rect 19716 89188 19740 89190
rect 19796 89188 19820 89190
rect 19876 89188 19882 89190
rect 19574 89168 19882 89188
rect 19574 88156 19882 88176
rect 19574 88154 19580 88156
rect 19636 88154 19660 88156
rect 19716 88154 19740 88156
rect 19796 88154 19820 88156
rect 19876 88154 19882 88156
rect 19636 88102 19638 88154
rect 19818 88102 19820 88154
rect 19574 88100 19580 88102
rect 19636 88100 19660 88102
rect 19716 88100 19740 88102
rect 19796 88100 19820 88102
rect 19876 88100 19882 88102
rect 19574 88080 19882 88100
rect 19574 87068 19882 87088
rect 19574 87066 19580 87068
rect 19636 87066 19660 87068
rect 19716 87066 19740 87068
rect 19796 87066 19820 87068
rect 19876 87066 19882 87068
rect 19636 87014 19638 87066
rect 19818 87014 19820 87066
rect 19574 87012 19580 87014
rect 19636 87012 19660 87014
rect 19716 87012 19740 87014
rect 19796 87012 19820 87014
rect 19876 87012 19882 87014
rect 19574 86992 19882 87012
rect 19574 85980 19882 86000
rect 19574 85978 19580 85980
rect 19636 85978 19660 85980
rect 19716 85978 19740 85980
rect 19796 85978 19820 85980
rect 19876 85978 19882 85980
rect 19636 85926 19638 85978
rect 19818 85926 19820 85978
rect 19574 85924 19580 85926
rect 19636 85924 19660 85926
rect 19716 85924 19740 85926
rect 19796 85924 19820 85926
rect 19876 85924 19882 85926
rect 19574 85904 19882 85924
rect 19574 84892 19882 84912
rect 19574 84890 19580 84892
rect 19636 84890 19660 84892
rect 19716 84890 19740 84892
rect 19796 84890 19820 84892
rect 19876 84890 19882 84892
rect 19636 84838 19638 84890
rect 19818 84838 19820 84890
rect 19574 84836 19580 84838
rect 19636 84836 19660 84838
rect 19716 84836 19740 84838
rect 19796 84836 19820 84838
rect 19876 84836 19882 84838
rect 19574 84816 19882 84836
rect 19574 83804 19882 83824
rect 19574 83802 19580 83804
rect 19636 83802 19660 83804
rect 19716 83802 19740 83804
rect 19796 83802 19820 83804
rect 19876 83802 19882 83804
rect 19636 83750 19638 83802
rect 19818 83750 19820 83802
rect 19574 83748 19580 83750
rect 19636 83748 19660 83750
rect 19716 83748 19740 83750
rect 19796 83748 19820 83750
rect 19876 83748 19882 83750
rect 19574 83728 19882 83748
rect 19574 82716 19882 82736
rect 19574 82714 19580 82716
rect 19636 82714 19660 82716
rect 19716 82714 19740 82716
rect 19796 82714 19820 82716
rect 19876 82714 19882 82716
rect 19636 82662 19638 82714
rect 19818 82662 19820 82714
rect 19574 82660 19580 82662
rect 19636 82660 19660 82662
rect 19716 82660 19740 82662
rect 19796 82660 19820 82662
rect 19876 82660 19882 82662
rect 19574 82640 19882 82660
rect 19574 81628 19882 81648
rect 19574 81626 19580 81628
rect 19636 81626 19660 81628
rect 19716 81626 19740 81628
rect 19796 81626 19820 81628
rect 19876 81626 19882 81628
rect 19636 81574 19638 81626
rect 19818 81574 19820 81626
rect 19574 81572 19580 81574
rect 19636 81572 19660 81574
rect 19716 81572 19740 81574
rect 19796 81572 19820 81574
rect 19876 81572 19882 81574
rect 19574 81552 19882 81572
rect 19574 80540 19882 80560
rect 19574 80538 19580 80540
rect 19636 80538 19660 80540
rect 19716 80538 19740 80540
rect 19796 80538 19820 80540
rect 19876 80538 19882 80540
rect 19636 80486 19638 80538
rect 19818 80486 19820 80538
rect 19574 80484 19580 80486
rect 19636 80484 19660 80486
rect 19716 80484 19740 80486
rect 19796 80484 19820 80486
rect 19876 80484 19882 80486
rect 19574 80464 19882 80484
rect 19574 79452 19882 79472
rect 19574 79450 19580 79452
rect 19636 79450 19660 79452
rect 19716 79450 19740 79452
rect 19796 79450 19820 79452
rect 19876 79450 19882 79452
rect 19636 79398 19638 79450
rect 19818 79398 19820 79450
rect 19574 79396 19580 79398
rect 19636 79396 19660 79398
rect 19716 79396 19740 79398
rect 19796 79396 19820 79398
rect 19876 79396 19882 79398
rect 19574 79376 19882 79396
rect 19574 78364 19882 78384
rect 19574 78362 19580 78364
rect 19636 78362 19660 78364
rect 19716 78362 19740 78364
rect 19796 78362 19820 78364
rect 19876 78362 19882 78364
rect 19636 78310 19638 78362
rect 19818 78310 19820 78362
rect 19574 78308 19580 78310
rect 19636 78308 19660 78310
rect 19716 78308 19740 78310
rect 19796 78308 19820 78310
rect 19876 78308 19882 78310
rect 19574 78288 19882 78308
rect 19574 77276 19882 77296
rect 19574 77274 19580 77276
rect 19636 77274 19660 77276
rect 19716 77274 19740 77276
rect 19796 77274 19820 77276
rect 19876 77274 19882 77276
rect 19636 77222 19638 77274
rect 19818 77222 19820 77274
rect 19574 77220 19580 77222
rect 19636 77220 19660 77222
rect 19716 77220 19740 77222
rect 19796 77220 19820 77222
rect 19876 77220 19882 77222
rect 19574 77200 19882 77220
rect 19574 76188 19882 76208
rect 19574 76186 19580 76188
rect 19636 76186 19660 76188
rect 19716 76186 19740 76188
rect 19796 76186 19820 76188
rect 19876 76186 19882 76188
rect 19636 76134 19638 76186
rect 19818 76134 19820 76186
rect 19574 76132 19580 76134
rect 19636 76132 19660 76134
rect 19716 76132 19740 76134
rect 19796 76132 19820 76134
rect 19876 76132 19882 76134
rect 19574 76112 19882 76132
rect 19574 75100 19882 75120
rect 19574 75098 19580 75100
rect 19636 75098 19660 75100
rect 19716 75098 19740 75100
rect 19796 75098 19820 75100
rect 19876 75098 19882 75100
rect 19636 75046 19638 75098
rect 19818 75046 19820 75098
rect 19574 75044 19580 75046
rect 19636 75044 19660 75046
rect 19716 75044 19740 75046
rect 19796 75044 19820 75046
rect 19876 75044 19882 75046
rect 19574 75024 19882 75044
rect 19574 74012 19882 74032
rect 19574 74010 19580 74012
rect 19636 74010 19660 74012
rect 19716 74010 19740 74012
rect 19796 74010 19820 74012
rect 19876 74010 19882 74012
rect 19636 73958 19638 74010
rect 19818 73958 19820 74010
rect 19574 73956 19580 73958
rect 19636 73956 19660 73958
rect 19716 73956 19740 73958
rect 19796 73956 19820 73958
rect 19876 73956 19882 73958
rect 19574 73936 19882 73956
rect 19574 72924 19882 72944
rect 19574 72922 19580 72924
rect 19636 72922 19660 72924
rect 19716 72922 19740 72924
rect 19796 72922 19820 72924
rect 19876 72922 19882 72924
rect 19636 72870 19638 72922
rect 19818 72870 19820 72922
rect 19574 72868 19580 72870
rect 19636 72868 19660 72870
rect 19716 72868 19740 72870
rect 19796 72868 19820 72870
rect 19876 72868 19882 72870
rect 19574 72848 19882 72868
rect 19574 71836 19882 71856
rect 19574 71834 19580 71836
rect 19636 71834 19660 71836
rect 19716 71834 19740 71836
rect 19796 71834 19820 71836
rect 19876 71834 19882 71836
rect 19636 71782 19638 71834
rect 19818 71782 19820 71834
rect 19574 71780 19580 71782
rect 19636 71780 19660 71782
rect 19716 71780 19740 71782
rect 19796 71780 19820 71782
rect 19876 71780 19882 71782
rect 19574 71760 19882 71780
rect 19574 70748 19882 70768
rect 19574 70746 19580 70748
rect 19636 70746 19660 70748
rect 19716 70746 19740 70748
rect 19796 70746 19820 70748
rect 19876 70746 19882 70748
rect 19636 70694 19638 70746
rect 19818 70694 19820 70746
rect 19574 70692 19580 70694
rect 19636 70692 19660 70694
rect 19716 70692 19740 70694
rect 19796 70692 19820 70694
rect 19876 70692 19882 70694
rect 19574 70672 19882 70692
rect 19574 69660 19882 69680
rect 19574 69658 19580 69660
rect 19636 69658 19660 69660
rect 19716 69658 19740 69660
rect 19796 69658 19820 69660
rect 19876 69658 19882 69660
rect 19636 69606 19638 69658
rect 19818 69606 19820 69658
rect 19574 69604 19580 69606
rect 19636 69604 19660 69606
rect 19716 69604 19740 69606
rect 19796 69604 19820 69606
rect 19876 69604 19882 69606
rect 19574 69584 19882 69604
rect 19574 68572 19882 68592
rect 19574 68570 19580 68572
rect 19636 68570 19660 68572
rect 19716 68570 19740 68572
rect 19796 68570 19820 68572
rect 19876 68570 19882 68572
rect 19636 68518 19638 68570
rect 19818 68518 19820 68570
rect 19574 68516 19580 68518
rect 19636 68516 19660 68518
rect 19716 68516 19740 68518
rect 19796 68516 19820 68518
rect 19876 68516 19882 68518
rect 19574 68496 19882 68516
rect 19574 67484 19882 67504
rect 19574 67482 19580 67484
rect 19636 67482 19660 67484
rect 19716 67482 19740 67484
rect 19796 67482 19820 67484
rect 19876 67482 19882 67484
rect 19636 67430 19638 67482
rect 19818 67430 19820 67482
rect 19574 67428 19580 67430
rect 19636 67428 19660 67430
rect 19716 67428 19740 67430
rect 19796 67428 19820 67430
rect 19876 67428 19882 67430
rect 19574 67408 19882 67428
rect 19574 66396 19882 66416
rect 19574 66394 19580 66396
rect 19636 66394 19660 66396
rect 19716 66394 19740 66396
rect 19796 66394 19820 66396
rect 19876 66394 19882 66396
rect 19636 66342 19638 66394
rect 19818 66342 19820 66394
rect 19574 66340 19580 66342
rect 19636 66340 19660 66342
rect 19716 66340 19740 66342
rect 19796 66340 19820 66342
rect 19876 66340 19882 66342
rect 19574 66320 19882 66340
rect 19574 65308 19882 65328
rect 19574 65306 19580 65308
rect 19636 65306 19660 65308
rect 19716 65306 19740 65308
rect 19796 65306 19820 65308
rect 19876 65306 19882 65308
rect 19636 65254 19638 65306
rect 19818 65254 19820 65306
rect 19574 65252 19580 65254
rect 19636 65252 19660 65254
rect 19716 65252 19740 65254
rect 19796 65252 19820 65254
rect 19876 65252 19882 65254
rect 19574 65232 19882 65252
rect 19574 64220 19882 64240
rect 19574 64218 19580 64220
rect 19636 64218 19660 64220
rect 19716 64218 19740 64220
rect 19796 64218 19820 64220
rect 19876 64218 19882 64220
rect 19636 64166 19638 64218
rect 19818 64166 19820 64218
rect 19574 64164 19580 64166
rect 19636 64164 19660 64166
rect 19716 64164 19740 64166
rect 19796 64164 19820 64166
rect 19876 64164 19882 64166
rect 19574 64144 19882 64164
rect 19574 63132 19882 63152
rect 19574 63130 19580 63132
rect 19636 63130 19660 63132
rect 19716 63130 19740 63132
rect 19796 63130 19820 63132
rect 19876 63130 19882 63132
rect 19636 63078 19638 63130
rect 19818 63078 19820 63130
rect 19574 63076 19580 63078
rect 19636 63076 19660 63078
rect 19716 63076 19740 63078
rect 19796 63076 19820 63078
rect 19876 63076 19882 63078
rect 19574 63056 19882 63076
rect 19574 62044 19882 62064
rect 19574 62042 19580 62044
rect 19636 62042 19660 62044
rect 19716 62042 19740 62044
rect 19796 62042 19820 62044
rect 19876 62042 19882 62044
rect 19636 61990 19638 62042
rect 19818 61990 19820 62042
rect 19574 61988 19580 61990
rect 19636 61988 19660 61990
rect 19716 61988 19740 61990
rect 19796 61988 19820 61990
rect 19876 61988 19882 61990
rect 19574 61968 19882 61988
rect 19432 61124 19484 61130
rect 19432 61066 19484 61072
rect 19574 60956 19882 60976
rect 19574 60954 19580 60956
rect 19636 60954 19660 60956
rect 19716 60954 19740 60956
rect 19796 60954 19820 60956
rect 19876 60954 19882 60956
rect 19636 60902 19638 60954
rect 19818 60902 19820 60954
rect 19574 60900 19580 60902
rect 19636 60900 19660 60902
rect 19716 60900 19740 60902
rect 19796 60900 19820 60902
rect 19876 60900 19882 60902
rect 19574 60880 19882 60900
rect 4214 60412 4522 60432
rect 4214 60410 4220 60412
rect 4276 60410 4300 60412
rect 4356 60410 4380 60412
rect 4436 60410 4460 60412
rect 4516 60410 4522 60412
rect 4276 60358 4278 60410
rect 4458 60358 4460 60410
rect 4214 60356 4220 60358
rect 4276 60356 4300 60358
rect 4356 60356 4380 60358
rect 4436 60356 4460 60358
rect 4516 60356 4522 60358
rect 4214 60336 4522 60356
rect 22664 60178 22692 117234
rect 22848 117162 22876 119326
rect 26422 119200 26478 120000
rect 30286 119200 30342 120000
rect 34150 119354 34206 120000
rect 37370 119354 37426 120000
rect 41234 119354 41290 120000
rect 45098 119354 45154 120000
rect 48962 119354 49018 120000
rect 52182 119354 52238 120000
rect 56046 119354 56102 120000
rect 34150 119326 34468 119354
rect 34150 119200 34206 119326
rect 26436 117298 26464 119200
rect 26424 117292 26476 117298
rect 26424 117234 26476 117240
rect 28264 117292 28316 117298
rect 28264 117234 28316 117240
rect 22836 117156 22888 117162
rect 22836 117098 22888 117104
rect 28276 114170 28304 117234
rect 30300 117178 30328 119200
rect 34440 117178 34468 119326
rect 37370 119326 37688 119354
rect 37370 119200 37426 119326
rect 34704 117292 34756 117298
rect 34704 117234 34756 117240
rect 36360 117292 36412 117298
rect 36360 117234 36412 117240
rect 30300 117162 30420 117178
rect 34440 117162 34560 117178
rect 30300 117156 30432 117162
rect 30300 117150 30380 117156
rect 34440 117156 34572 117162
rect 34440 117150 34520 117156
rect 30380 117098 30432 117104
rect 34520 117098 34572 117104
rect 34716 116822 34744 117234
rect 35808 117224 35860 117230
rect 35808 117166 35860 117172
rect 34934 116988 35242 117008
rect 34934 116986 34940 116988
rect 34996 116986 35020 116988
rect 35076 116986 35100 116988
rect 35156 116986 35180 116988
rect 35236 116986 35242 116988
rect 34996 116934 34998 116986
rect 35178 116934 35180 116986
rect 34934 116932 34940 116934
rect 34996 116932 35020 116934
rect 35076 116932 35100 116934
rect 35156 116932 35180 116934
rect 35236 116932 35242 116934
rect 34934 116912 35242 116932
rect 34704 116816 34756 116822
rect 34704 116758 34756 116764
rect 34934 115900 35242 115920
rect 34934 115898 34940 115900
rect 34996 115898 35020 115900
rect 35076 115898 35100 115900
rect 35156 115898 35180 115900
rect 35236 115898 35242 115900
rect 34996 115846 34998 115898
rect 35178 115846 35180 115898
rect 34934 115844 34940 115846
rect 34996 115844 35020 115846
rect 35076 115844 35100 115846
rect 35156 115844 35180 115846
rect 35236 115844 35242 115846
rect 34934 115824 35242 115844
rect 34934 114812 35242 114832
rect 34934 114810 34940 114812
rect 34996 114810 35020 114812
rect 35076 114810 35100 114812
rect 35156 114810 35180 114812
rect 35236 114810 35242 114812
rect 34996 114758 34998 114810
rect 35178 114758 35180 114810
rect 34934 114756 34940 114758
rect 34996 114756 35020 114758
rect 35076 114756 35100 114758
rect 35156 114756 35180 114758
rect 35236 114756 35242 114758
rect 34934 114736 35242 114756
rect 28264 114164 28316 114170
rect 28264 114106 28316 114112
rect 34934 113724 35242 113744
rect 34934 113722 34940 113724
rect 34996 113722 35020 113724
rect 35076 113722 35100 113724
rect 35156 113722 35180 113724
rect 35236 113722 35242 113724
rect 34996 113670 34998 113722
rect 35178 113670 35180 113722
rect 34934 113668 34940 113670
rect 34996 113668 35020 113670
rect 35076 113668 35100 113670
rect 35156 113668 35180 113670
rect 35236 113668 35242 113670
rect 34934 113648 35242 113668
rect 34934 112636 35242 112656
rect 34934 112634 34940 112636
rect 34996 112634 35020 112636
rect 35076 112634 35100 112636
rect 35156 112634 35180 112636
rect 35236 112634 35242 112636
rect 34996 112582 34998 112634
rect 35178 112582 35180 112634
rect 34934 112580 34940 112582
rect 34996 112580 35020 112582
rect 35076 112580 35100 112582
rect 35156 112580 35180 112582
rect 35236 112580 35242 112582
rect 34934 112560 35242 112580
rect 34934 111548 35242 111568
rect 34934 111546 34940 111548
rect 34996 111546 35020 111548
rect 35076 111546 35100 111548
rect 35156 111546 35180 111548
rect 35236 111546 35242 111548
rect 34996 111494 34998 111546
rect 35178 111494 35180 111546
rect 34934 111492 34940 111494
rect 34996 111492 35020 111494
rect 35076 111492 35100 111494
rect 35156 111492 35180 111494
rect 35236 111492 35242 111494
rect 34934 111472 35242 111492
rect 34934 110460 35242 110480
rect 34934 110458 34940 110460
rect 34996 110458 35020 110460
rect 35076 110458 35100 110460
rect 35156 110458 35180 110460
rect 35236 110458 35242 110460
rect 34996 110406 34998 110458
rect 35178 110406 35180 110458
rect 34934 110404 34940 110406
rect 34996 110404 35020 110406
rect 35076 110404 35100 110406
rect 35156 110404 35180 110406
rect 35236 110404 35242 110406
rect 34934 110384 35242 110404
rect 34934 109372 35242 109392
rect 34934 109370 34940 109372
rect 34996 109370 35020 109372
rect 35076 109370 35100 109372
rect 35156 109370 35180 109372
rect 35236 109370 35242 109372
rect 34996 109318 34998 109370
rect 35178 109318 35180 109370
rect 34934 109316 34940 109318
rect 34996 109316 35020 109318
rect 35076 109316 35100 109318
rect 35156 109316 35180 109318
rect 35236 109316 35242 109318
rect 34934 109296 35242 109316
rect 34934 108284 35242 108304
rect 34934 108282 34940 108284
rect 34996 108282 35020 108284
rect 35076 108282 35100 108284
rect 35156 108282 35180 108284
rect 35236 108282 35242 108284
rect 34996 108230 34998 108282
rect 35178 108230 35180 108282
rect 34934 108228 34940 108230
rect 34996 108228 35020 108230
rect 35076 108228 35100 108230
rect 35156 108228 35180 108230
rect 35236 108228 35242 108230
rect 34934 108208 35242 108228
rect 34934 107196 35242 107216
rect 34934 107194 34940 107196
rect 34996 107194 35020 107196
rect 35076 107194 35100 107196
rect 35156 107194 35180 107196
rect 35236 107194 35242 107196
rect 34996 107142 34998 107194
rect 35178 107142 35180 107194
rect 34934 107140 34940 107142
rect 34996 107140 35020 107142
rect 35076 107140 35100 107142
rect 35156 107140 35180 107142
rect 35236 107140 35242 107142
rect 34934 107120 35242 107140
rect 34934 106108 35242 106128
rect 34934 106106 34940 106108
rect 34996 106106 35020 106108
rect 35076 106106 35100 106108
rect 35156 106106 35180 106108
rect 35236 106106 35242 106108
rect 34996 106054 34998 106106
rect 35178 106054 35180 106106
rect 34934 106052 34940 106054
rect 34996 106052 35020 106054
rect 35076 106052 35100 106054
rect 35156 106052 35180 106054
rect 35236 106052 35242 106054
rect 34934 106032 35242 106052
rect 34934 105020 35242 105040
rect 34934 105018 34940 105020
rect 34996 105018 35020 105020
rect 35076 105018 35100 105020
rect 35156 105018 35180 105020
rect 35236 105018 35242 105020
rect 34996 104966 34998 105018
rect 35178 104966 35180 105018
rect 34934 104964 34940 104966
rect 34996 104964 35020 104966
rect 35076 104964 35100 104966
rect 35156 104964 35180 104966
rect 35236 104964 35242 104966
rect 34934 104944 35242 104964
rect 34934 103932 35242 103952
rect 34934 103930 34940 103932
rect 34996 103930 35020 103932
rect 35076 103930 35100 103932
rect 35156 103930 35180 103932
rect 35236 103930 35242 103932
rect 34996 103878 34998 103930
rect 35178 103878 35180 103930
rect 34934 103876 34940 103878
rect 34996 103876 35020 103878
rect 35076 103876 35100 103878
rect 35156 103876 35180 103878
rect 35236 103876 35242 103878
rect 34934 103856 35242 103876
rect 34934 102844 35242 102864
rect 34934 102842 34940 102844
rect 34996 102842 35020 102844
rect 35076 102842 35100 102844
rect 35156 102842 35180 102844
rect 35236 102842 35242 102844
rect 34996 102790 34998 102842
rect 35178 102790 35180 102842
rect 34934 102788 34940 102790
rect 34996 102788 35020 102790
rect 35076 102788 35100 102790
rect 35156 102788 35180 102790
rect 35236 102788 35242 102790
rect 34934 102768 35242 102788
rect 34934 101756 35242 101776
rect 34934 101754 34940 101756
rect 34996 101754 35020 101756
rect 35076 101754 35100 101756
rect 35156 101754 35180 101756
rect 35236 101754 35242 101756
rect 34996 101702 34998 101754
rect 35178 101702 35180 101754
rect 34934 101700 34940 101702
rect 34996 101700 35020 101702
rect 35076 101700 35100 101702
rect 35156 101700 35180 101702
rect 35236 101700 35242 101702
rect 34934 101680 35242 101700
rect 34934 100668 35242 100688
rect 34934 100666 34940 100668
rect 34996 100666 35020 100668
rect 35076 100666 35100 100668
rect 35156 100666 35180 100668
rect 35236 100666 35242 100668
rect 34996 100614 34998 100666
rect 35178 100614 35180 100666
rect 34934 100612 34940 100614
rect 34996 100612 35020 100614
rect 35076 100612 35100 100614
rect 35156 100612 35180 100614
rect 35236 100612 35242 100614
rect 34934 100592 35242 100612
rect 34934 99580 35242 99600
rect 34934 99578 34940 99580
rect 34996 99578 35020 99580
rect 35076 99578 35100 99580
rect 35156 99578 35180 99580
rect 35236 99578 35242 99580
rect 34996 99526 34998 99578
rect 35178 99526 35180 99578
rect 34934 99524 34940 99526
rect 34996 99524 35020 99526
rect 35076 99524 35100 99526
rect 35156 99524 35180 99526
rect 35236 99524 35242 99526
rect 34934 99504 35242 99524
rect 34934 98492 35242 98512
rect 34934 98490 34940 98492
rect 34996 98490 35020 98492
rect 35076 98490 35100 98492
rect 35156 98490 35180 98492
rect 35236 98490 35242 98492
rect 34996 98438 34998 98490
rect 35178 98438 35180 98490
rect 34934 98436 34940 98438
rect 34996 98436 35020 98438
rect 35076 98436 35100 98438
rect 35156 98436 35180 98438
rect 35236 98436 35242 98438
rect 34934 98416 35242 98436
rect 34934 97404 35242 97424
rect 34934 97402 34940 97404
rect 34996 97402 35020 97404
rect 35076 97402 35100 97404
rect 35156 97402 35180 97404
rect 35236 97402 35242 97404
rect 34996 97350 34998 97402
rect 35178 97350 35180 97402
rect 34934 97348 34940 97350
rect 34996 97348 35020 97350
rect 35076 97348 35100 97350
rect 35156 97348 35180 97350
rect 35236 97348 35242 97350
rect 34934 97328 35242 97348
rect 34934 96316 35242 96336
rect 34934 96314 34940 96316
rect 34996 96314 35020 96316
rect 35076 96314 35100 96316
rect 35156 96314 35180 96316
rect 35236 96314 35242 96316
rect 34996 96262 34998 96314
rect 35178 96262 35180 96314
rect 34934 96260 34940 96262
rect 34996 96260 35020 96262
rect 35076 96260 35100 96262
rect 35156 96260 35180 96262
rect 35236 96260 35242 96262
rect 34934 96240 35242 96260
rect 34934 95228 35242 95248
rect 34934 95226 34940 95228
rect 34996 95226 35020 95228
rect 35076 95226 35100 95228
rect 35156 95226 35180 95228
rect 35236 95226 35242 95228
rect 34996 95174 34998 95226
rect 35178 95174 35180 95226
rect 34934 95172 34940 95174
rect 34996 95172 35020 95174
rect 35076 95172 35100 95174
rect 35156 95172 35180 95174
rect 35236 95172 35242 95174
rect 34934 95152 35242 95172
rect 34934 94140 35242 94160
rect 34934 94138 34940 94140
rect 34996 94138 35020 94140
rect 35076 94138 35100 94140
rect 35156 94138 35180 94140
rect 35236 94138 35242 94140
rect 34996 94086 34998 94138
rect 35178 94086 35180 94138
rect 34934 94084 34940 94086
rect 34996 94084 35020 94086
rect 35076 94084 35100 94086
rect 35156 94084 35180 94086
rect 35236 94084 35242 94086
rect 34934 94064 35242 94084
rect 34934 93052 35242 93072
rect 34934 93050 34940 93052
rect 34996 93050 35020 93052
rect 35076 93050 35100 93052
rect 35156 93050 35180 93052
rect 35236 93050 35242 93052
rect 34996 92998 34998 93050
rect 35178 92998 35180 93050
rect 34934 92996 34940 92998
rect 34996 92996 35020 92998
rect 35076 92996 35100 92998
rect 35156 92996 35180 92998
rect 35236 92996 35242 92998
rect 34934 92976 35242 92996
rect 34934 91964 35242 91984
rect 34934 91962 34940 91964
rect 34996 91962 35020 91964
rect 35076 91962 35100 91964
rect 35156 91962 35180 91964
rect 35236 91962 35242 91964
rect 34996 91910 34998 91962
rect 35178 91910 35180 91962
rect 34934 91908 34940 91910
rect 34996 91908 35020 91910
rect 35076 91908 35100 91910
rect 35156 91908 35180 91910
rect 35236 91908 35242 91910
rect 34934 91888 35242 91908
rect 34934 90876 35242 90896
rect 34934 90874 34940 90876
rect 34996 90874 35020 90876
rect 35076 90874 35100 90876
rect 35156 90874 35180 90876
rect 35236 90874 35242 90876
rect 34996 90822 34998 90874
rect 35178 90822 35180 90874
rect 34934 90820 34940 90822
rect 34996 90820 35020 90822
rect 35076 90820 35100 90822
rect 35156 90820 35180 90822
rect 35236 90820 35242 90822
rect 34934 90800 35242 90820
rect 34934 89788 35242 89808
rect 34934 89786 34940 89788
rect 34996 89786 35020 89788
rect 35076 89786 35100 89788
rect 35156 89786 35180 89788
rect 35236 89786 35242 89788
rect 34996 89734 34998 89786
rect 35178 89734 35180 89786
rect 34934 89732 34940 89734
rect 34996 89732 35020 89734
rect 35076 89732 35100 89734
rect 35156 89732 35180 89734
rect 35236 89732 35242 89734
rect 34934 89712 35242 89732
rect 34934 88700 35242 88720
rect 34934 88698 34940 88700
rect 34996 88698 35020 88700
rect 35076 88698 35100 88700
rect 35156 88698 35180 88700
rect 35236 88698 35242 88700
rect 34996 88646 34998 88698
rect 35178 88646 35180 88698
rect 34934 88644 34940 88646
rect 34996 88644 35020 88646
rect 35076 88644 35100 88646
rect 35156 88644 35180 88646
rect 35236 88644 35242 88646
rect 34934 88624 35242 88644
rect 34934 87612 35242 87632
rect 34934 87610 34940 87612
rect 34996 87610 35020 87612
rect 35076 87610 35100 87612
rect 35156 87610 35180 87612
rect 35236 87610 35242 87612
rect 34996 87558 34998 87610
rect 35178 87558 35180 87610
rect 34934 87556 34940 87558
rect 34996 87556 35020 87558
rect 35076 87556 35100 87558
rect 35156 87556 35180 87558
rect 35236 87556 35242 87558
rect 34934 87536 35242 87556
rect 34934 86524 35242 86544
rect 34934 86522 34940 86524
rect 34996 86522 35020 86524
rect 35076 86522 35100 86524
rect 35156 86522 35180 86524
rect 35236 86522 35242 86524
rect 34996 86470 34998 86522
rect 35178 86470 35180 86522
rect 34934 86468 34940 86470
rect 34996 86468 35020 86470
rect 35076 86468 35100 86470
rect 35156 86468 35180 86470
rect 35236 86468 35242 86470
rect 34934 86448 35242 86468
rect 34934 85436 35242 85456
rect 34934 85434 34940 85436
rect 34996 85434 35020 85436
rect 35076 85434 35100 85436
rect 35156 85434 35180 85436
rect 35236 85434 35242 85436
rect 34996 85382 34998 85434
rect 35178 85382 35180 85434
rect 34934 85380 34940 85382
rect 34996 85380 35020 85382
rect 35076 85380 35100 85382
rect 35156 85380 35180 85382
rect 35236 85380 35242 85382
rect 34934 85360 35242 85380
rect 34934 84348 35242 84368
rect 34934 84346 34940 84348
rect 34996 84346 35020 84348
rect 35076 84346 35100 84348
rect 35156 84346 35180 84348
rect 35236 84346 35242 84348
rect 34996 84294 34998 84346
rect 35178 84294 35180 84346
rect 34934 84292 34940 84294
rect 34996 84292 35020 84294
rect 35076 84292 35100 84294
rect 35156 84292 35180 84294
rect 35236 84292 35242 84294
rect 34934 84272 35242 84292
rect 34934 83260 35242 83280
rect 34934 83258 34940 83260
rect 34996 83258 35020 83260
rect 35076 83258 35100 83260
rect 35156 83258 35180 83260
rect 35236 83258 35242 83260
rect 34996 83206 34998 83258
rect 35178 83206 35180 83258
rect 34934 83204 34940 83206
rect 34996 83204 35020 83206
rect 35076 83204 35100 83206
rect 35156 83204 35180 83206
rect 35236 83204 35242 83206
rect 34934 83184 35242 83204
rect 34934 82172 35242 82192
rect 34934 82170 34940 82172
rect 34996 82170 35020 82172
rect 35076 82170 35100 82172
rect 35156 82170 35180 82172
rect 35236 82170 35242 82172
rect 34996 82118 34998 82170
rect 35178 82118 35180 82170
rect 34934 82116 34940 82118
rect 34996 82116 35020 82118
rect 35076 82116 35100 82118
rect 35156 82116 35180 82118
rect 35236 82116 35242 82118
rect 34934 82096 35242 82116
rect 34934 81084 35242 81104
rect 34934 81082 34940 81084
rect 34996 81082 35020 81084
rect 35076 81082 35100 81084
rect 35156 81082 35180 81084
rect 35236 81082 35242 81084
rect 34996 81030 34998 81082
rect 35178 81030 35180 81082
rect 34934 81028 34940 81030
rect 34996 81028 35020 81030
rect 35076 81028 35100 81030
rect 35156 81028 35180 81030
rect 35236 81028 35242 81030
rect 34934 81008 35242 81028
rect 34934 79996 35242 80016
rect 34934 79994 34940 79996
rect 34996 79994 35020 79996
rect 35076 79994 35100 79996
rect 35156 79994 35180 79996
rect 35236 79994 35242 79996
rect 34996 79942 34998 79994
rect 35178 79942 35180 79994
rect 34934 79940 34940 79942
rect 34996 79940 35020 79942
rect 35076 79940 35100 79942
rect 35156 79940 35180 79942
rect 35236 79940 35242 79942
rect 34934 79920 35242 79940
rect 34934 78908 35242 78928
rect 34934 78906 34940 78908
rect 34996 78906 35020 78908
rect 35076 78906 35100 78908
rect 35156 78906 35180 78908
rect 35236 78906 35242 78908
rect 34996 78854 34998 78906
rect 35178 78854 35180 78906
rect 34934 78852 34940 78854
rect 34996 78852 35020 78854
rect 35076 78852 35100 78854
rect 35156 78852 35180 78854
rect 35236 78852 35242 78854
rect 34934 78832 35242 78852
rect 34934 77820 35242 77840
rect 34934 77818 34940 77820
rect 34996 77818 35020 77820
rect 35076 77818 35100 77820
rect 35156 77818 35180 77820
rect 35236 77818 35242 77820
rect 34996 77766 34998 77818
rect 35178 77766 35180 77818
rect 34934 77764 34940 77766
rect 34996 77764 35020 77766
rect 35076 77764 35100 77766
rect 35156 77764 35180 77766
rect 35236 77764 35242 77766
rect 34934 77744 35242 77764
rect 34934 76732 35242 76752
rect 34934 76730 34940 76732
rect 34996 76730 35020 76732
rect 35076 76730 35100 76732
rect 35156 76730 35180 76732
rect 35236 76730 35242 76732
rect 34996 76678 34998 76730
rect 35178 76678 35180 76730
rect 34934 76676 34940 76678
rect 34996 76676 35020 76678
rect 35076 76676 35100 76678
rect 35156 76676 35180 76678
rect 35236 76676 35242 76678
rect 34934 76656 35242 76676
rect 34934 75644 35242 75664
rect 34934 75642 34940 75644
rect 34996 75642 35020 75644
rect 35076 75642 35100 75644
rect 35156 75642 35180 75644
rect 35236 75642 35242 75644
rect 34996 75590 34998 75642
rect 35178 75590 35180 75642
rect 34934 75588 34940 75590
rect 34996 75588 35020 75590
rect 35076 75588 35100 75590
rect 35156 75588 35180 75590
rect 35236 75588 35242 75590
rect 34934 75568 35242 75588
rect 34934 74556 35242 74576
rect 34934 74554 34940 74556
rect 34996 74554 35020 74556
rect 35076 74554 35100 74556
rect 35156 74554 35180 74556
rect 35236 74554 35242 74556
rect 34996 74502 34998 74554
rect 35178 74502 35180 74554
rect 34934 74500 34940 74502
rect 34996 74500 35020 74502
rect 35076 74500 35100 74502
rect 35156 74500 35180 74502
rect 35236 74500 35242 74502
rect 34934 74480 35242 74500
rect 34934 73468 35242 73488
rect 34934 73466 34940 73468
rect 34996 73466 35020 73468
rect 35076 73466 35100 73468
rect 35156 73466 35180 73468
rect 35236 73466 35242 73468
rect 34996 73414 34998 73466
rect 35178 73414 35180 73466
rect 34934 73412 34940 73414
rect 34996 73412 35020 73414
rect 35076 73412 35100 73414
rect 35156 73412 35180 73414
rect 35236 73412 35242 73414
rect 34934 73392 35242 73412
rect 34934 72380 35242 72400
rect 34934 72378 34940 72380
rect 34996 72378 35020 72380
rect 35076 72378 35100 72380
rect 35156 72378 35180 72380
rect 35236 72378 35242 72380
rect 34996 72326 34998 72378
rect 35178 72326 35180 72378
rect 34934 72324 34940 72326
rect 34996 72324 35020 72326
rect 35076 72324 35100 72326
rect 35156 72324 35180 72326
rect 35236 72324 35242 72326
rect 34934 72304 35242 72324
rect 34934 71292 35242 71312
rect 34934 71290 34940 71292
rect 34996 71290 35020 71292
rect 35076 71290 35100 71292
rect 35156 71290 35180 71292
rect 35236 71290 35242 71292
rect 34996 71238 34998 71290
rect 35178 71238 35180 71290
rect 34934 71236 34940 71238
rect 34996 71236 35020 71238
rect 35076 71236 35100 71238
rect 35156 71236 35180 71238
rect 35236 71236 35242 71238
rect 34934 71216 35242 71236
rect 34934 70204 35242 70224
rect 34934 70202 34940 70204
rect 34996 70202 35020 70204
rect 35076 70202 35100 70204
rect 35156 70202 35180 70204
rect 35236 70202 35242 70204
rect 34996 70150 34998 70202
rect 35178 70150 35180 70202
rect 34934 70148 34940 70150
rect 34996 70148 35020 70150
rect 35076 70148 35100 70150
rect 35156 70148 35180 70150
rect 35236 70148 35242 70150
rect 34934 70128 35242 70148
rect 34934 69116 35242 69136
rect 34934 69114 34940 69116
rect 34996 69114 35020 69116
rect 35076 69114 35100 69116
rect 35156 69114 35180 69116
rect 35236 69114 35242 69116
rect 34996 69062 34998 69114
rect 35178 69062 35180 69114
rect 34934 69060 34940 69062
rect 34996 69060 35020 69062
rect 35076 69060 35100 69062
rect 35156 69060 35180 69062
rect 35236 69060 35242 69062
rect 34934 69040 35242 69060
rect 34934 68028 35242 68048
rect 34934 68026 34940 68028
rect 34996 68026 35020 68028
rect 35076 68026 35100 68028
rect 35156 68026 35180 68028
rect 35236 68026 35242 68028
rect 34996 67974 34998 68026
rect 35178 67974 35180 68026
rect 34934 67972 34940 67974
rect 34996 67972 35020 67974
rect 35076 67972 35100 67974
rect 35156 67972 35180 67974
rect 35236 67972 35242 67974
rect 34934 67952 35242 67972
rect 34934 66940 35242 66960
rect 34934 66938 34940 66940
rect 34996 66938 35020 66940
rect 35076 66938 35100 66940
rect 35156 66938 35180 66940
rect 35236 66938 35242 66940
rect 34996 66886 34998 66938
rect 35178 66886 35180 66938
rect 34934 66884 34940 66886
rect 34996 66884 35020 66886
rect 35076 66884 35100 66886
rect 35156 66884 35180 66886
rect 35236 66884 35242 66886
rect 34934 66864 35242 66884
rect 34934 65852 35242 65872
rect 34934 65850 34940 65852
rect 34996 65850 35020 65852
rect 35076 65850 35100 65852
rect 35156 65850 35180 65852
rect 35236 65850 35242 65852
rect 34996 65798 34998 65850
rect 35178 65798 35180 65850
rect 34934 65796 34940 65798
rect 34996 65796 35020 65798
rect 35076 65796 35100 65798
rect 35156 65796 35180 65798
rect 35236 65796 35242 65798
rect 34934 65776 35242 65796
rect 34934 64764 35242 64784
rect 34934 64762 34940 64764
rect 34996 64762 35020 64764
rect 35076 64762 35100 64764
rect 35156 64762 35180 64764
rect 35236 64762 35242 64764
rect 34996 64710 34998 64762
rect 35178 64710 35180 64762
rect 34934 64708 34940 64710
rect 34996 64708 35020 64710
rect 35076 64708 35100 64710
rect 35156 64708 35180 64710
rect 35236 64708 35242 64710
rect 34934 64688 35242 64708
rect 34934 63676 35242 63696
rect 34934 63674 34940 63676
rect 34996 63674 35020 63676
rect 35076 63674 35100 63676
rect 35156 63674 35180 63676
rect 35236 63674 35242 63676
rect 34996 63622 34998 63674
rect 35178 63622 35180 63674
rect 34934 63620 34940 63622
rect 34996 63620 35020 63622
rect 35076 63620 35100 63622
rect 35156 63620 35180 63622
rect 35236 63620 35242 63622
rect 34934 63600 35242 63620
rect 34934 62588 35242 62608
rect 34934 62586 34940 62588
rect 34996 62586 35020 62588
rect 35076 62586 35100 62588
rect 35156 62586 35180 62588
rect 35236 62586 35242 62588
rect 34996 62534 34998 62586
rect 35178 62534 35180 62586
rect 34934 62532 34940 62534
rect 34996 62532 35020 62534
rect 35076 62532 35100 62534
rect 35156 62532 35180 62534
rect 35236 62532 35242 62534
rect 34934 62512 35242 62532
rect 34934 61500 35242 61520
rect 34934 61498 34940 61500
rect 34996 61498 35020 61500
rect 35076 61498 35100 61500
rect 35156 61498 35180 61500
rect 35236 61498 35242 61500
rect 34996 61446 34998 61498
rect 35178 61446 35180 61498
rect 34934 61444 34940 61446
rect 34996 61444 35020 61446
rect 35076 61444 35100 61446
rect 35156 61444 35180 61446
rect 35236 61444 35242 61446
rect 34934 61424 35242 61444
rect 34934 60412 35242 60432
rect 34934 60410 34940 60412
rect 34996 60410 35020 60412
rect 35076 60410 35100 60412
rect 35156 60410 35180 60412
rect 35236 60410 35242 60412
rect 34996 60358 34998 60410
rect 35178 60358 35180 60410
rect 34934 60356 34940 60358
rect 34996 60356 35020 60358
rect 35076 60356 35100 60358
rect 35156 60356 35180 60358
rect 35236 60356 35242 60358
rect 34934 60336 35242 60356
rect 35820 60314 35848 117166
rect 36372 60314 36400 117234
rect 37660 117162 37688 119326
rect 41234 119326 41368 119354
rect 41234 119200 41290 119326
rect 40684 117292 40736 117298
rect 40684 117234 40736 117240
rect 37464 117156 37516 117162
rect 37464 117098 37516 117104
rect 37648 117156 37700 117162
rect 37648 117098 37700 117104
rect 37476 116210 37504 117098
rect 40040 116748 40092 116754
rect 40040 116690 40092 116696
rect 37464 116204 37516 116210
rect 37464 116146 37516 116152
rect 40052 109274 40080 116690
rect 40040 109268 40092 109274
rect 40040 109210 40092 109216
rect 39856 109064 39908 109070
rect 39856 109006 39908 109012
rect 39868 101318 39896 109006
rect 39856 101312 39908 101318
rect 39856 101254 39908 101260
rect 40316 95940 40368 95946
rect 40316 95882 40368 95888
rect 39948 89004 40000 89010
rect 39948 88946 40000 88952
rect 39960 79014 39988 88946
rect 40328 87174 40356 95882
rect 40316 87168 40368 87174
rect 40316 87110 40368 87116
rect 39948 79008 40000 79014
rect 39948 78950 40000 78956
rect 40696 65618 40724 117234
rect 41340 117212 41368 119326
rect 45098 119326 45416 119354
rect 45098 119200 45154 119326
rect 45192 117292 45244 117298
rect 45192 117234 45244 117240
rect 41340 117184 41460 117212
rect 41432 117094 41460 117184
rect 41420 117088 41472 117094
rect 41420 117030 41472 117036
rect 40776 116884 40828 116890
rect 40776 116826 40828 116832
rect 41420 116884 41472 116890
rect 41420 116826 41472 116832
rect 40788 116346 40816 116826
rect 40776 116340 40828 116346
rect 40776 116282 40828 116288
rect 41432 92410 41460 116826
rect 41420 92404 41472 92410
rect 41420 92346 41472 92352
rect 41052 92268 41104 92274
rect 41052 92210 41104 92216
rect 41064 90030 41092 92210
rect 41052 90024 41104 90030
rect 41052 89966 41104 89972
rect 40684 65612 40736 65618
rect 40684 65554 40736 65560
rect 39856 65544 39908 65550
rect 39856 65486 39908 65492
rect 39488 64456 39540 64462
rect 39488 64398 39540 64404
rect 39500 63986 39528 64398
rect 39488 63980 39540 63986
rect 39488 63922 39540 63928
rect 39488 63776 39540 63782
rect 39488 63718 39540 63724
rect 38292 63368 38344 63374
rect 38292 63310 38344 63316
rect 38304 60314 38332 63310
rect 38844 60716 38896 60722
rect 38844 60658 38896 60664
rect 35808 60308 35860 60314
rect 35808 60250 35860 60256
rect 36360 60308 36412 60314
rect 36360 60250 36412 60256
rect 38292 60308 38344 60314
rect 38292 60250 38344 60256
rect 22652 60172 22704 60178
rect 22652 60114 22704 60120
rect 35820 60042 35848 60250
rect 19984 60036 20036 60042
rect 19984 59978 20036 59984
rect 35808 60036 35860 60042
rect 35808 59978 35860 59984
rect 36268 60036 36320 60042
rect 36268 59978 36320 59984
rect 19574 59868 19882 59888
rect 19574 59866 19580 59868
rect 19636 59866 19660 59868
rect 19716 59866 19740 59868
rect 19796 59866 19820 59868
rect 19876 59866 19882 59868
rect 19636 59814 19638 59866
rect 19818 59814 19820 59866
rect 19574 59812 19580 59814
rect 19636 59812 19660 59814
rect 19716 59812 19740 59814
rect 19796 59812 19820 59814
rect 19876 59812 19882 59814
rect 19574 59792 19882 59812
rect 4620 59764 4672 59770
rect 4620 59706 4672 59712
rect 4214 59324 4522 59344
rect 4214 59322 4220 59324
rect 4276 59322 4300 59324
rect 4356 59322 4380 59324
rect 4436 59322 4460 59324
rect 4516 59322 4522 59324
rect 4276 59270 4278 59322
rect 4458 59270 4460 59322
rect 4214 59268 4220 59270
rect 4276 59268 4300 59270
rect 4356 59268 4380 59270
rect 4436 59268 4460 59270
rect 4516 59268 4522 59270
rect 4214 59248 4522 59268
rect 4214 58236 4522 58256
rect 4214 58234 4220 58236
rect 4276 58234 4300 58236
rect 4356 58234 4380 58236
rect 4436 58234 4460 58236
rect 4516 58234 4522 58236
rect 4276 58182 4278 58234
rect 4458 58182 4460 58234
rect 4214 58180 4220 58182
rect 4276 58180 4300 58182
rect 4356 58180 4380 58182
rect 4436 58180 4460 58182
rect 4516 58180 4522 58182
rect 4214 58160 4522 58180
rect 4214 57148 4522 57168
rect 4214 57146 4220 57148
rect 4276 57146 4300 57148
rect 4356 57146 4380 57148
rect 4436 57146 4460 57148
rect 4516 57146 4522 57148
rect 4276 57094 4278 57146
rect 4458 57094 4460 57146
rect 4214 57092 4220 57094
rect 4276 57092 4300 57094
rect 4356 57092 4380 57094
rect 4436 57092 4460 57094
rect 4516 57092 4522 57094
rect 4214 57072 4522 57092
rect 4214 56060 4522 56080
rect 4214 56058 4220 56060
rect 4276 56058 4300 56060
rect 4356 56058 4380 56060
rect 4436 56058 4460 56060
rect 4516 56058 4522 56060
rect 4276 56006 4278 56058
rect 4458 56006 4460 56058
rect 4214 56004 4220 56006
rect 4276 56004 4300 56006
rect 4356 56004 4380 56006
rect 4436 56004 4460 56006
rect 4516 56004 4522 56006
rect 4214 55984 4522 56004
rect 4214 54972 4522 54992
rect 4214 54970 4220 54972
rect 4276 54970 4300 54972
rect 4356 54970 4380 54972
rect 4436 54970 4460 54972
rect 4516 54970 4522 54972
rect 4276 54918 4278 54970
rect 4458 54918 4460 54970
rect 4214 54916 4220 54918
rect 4276 54916 4300 54918
rect 4356 54916 4380 54918
rect 4436 54916 4460 54918
rect 4516 54916 4522 54918
rect 4214 54896 4522 54916
rect 4214 53884 4522 53904
rect 4214 53882 4220 53884
rect 4276 53882 4300 53884
rect 4356 53882 4380 53884
rect 4436 53882 4460 53884
rect 4516 53882 4522 53884
rect 4276 53830 4278 53882
rect 4458 53830 4460 53882
rect 4214 53828 4220 53830
rect 4276 53828 4300 53830
rect 4356 53828 4380 53830
rect 4436 53828 4460 53830
rect 4516 53828 4522 53830
rect 4214 53808 4522 53828
rect 4214 52796 4522 52816
rect 4214 52794 4220 52796
rect 4276 52794 4300 52796
rect 4356 52794 4380 52796
rect 4436 52794 4460 52796
rect 4516 52794 4522 52796
rect 4276 52742 4278 52794
rect 4458 52742 4460 52794
rect 4214 52740 4220 52742
rect 4276 52740 4300 52742
rect 4356 52740 4380 52742
rect 4436 52740 4460 52742
rect 4516 52740 4522 52742
rect 4214 52720 4522 52740
rect 4214 51708 4522 51728
rect 4214 51706 4220 51708
rect 4276 51706 4300 51708
rect 4356 51706 4380 51708
rect 4436 51706 4460 51708
rect 4516 51706 4522 51708
rect 4276 51654 4278 51706
rect 4458 51654 4460 51706
rect 4214 51652 4220 51654
rect 4276 51652 4300 51654
rect 4356 51652 4380 51654
rect 4436 51652 4460 51654
rect 4516 51652 4522 51654
rect 4214 51632 4522 51652
rect 4214 50620 4522 50640
rect 4214 50618 4220 50620
rect 4276 50618 4300 50620
rect 4356 50618 4380 50620
rect 4436 50618 4460 50620
rect 4516 50618 4522 50620
rect 4276 50566 4278 50618
rect 4458 50566 4460 50618
rect 4214 50564 4220 50566
rect 4276 50564 4300 50566
rect 4356 50564 4380 50566
rect 4436 50564 4460 50566
rect 4516 50564 4522 50566
rect 4214 50544 4522 50564
rect 4214 49532 4522 49552
rect 4214 49530 4220 49532
rect 4276 49530 4300 49532
rect 4356 49530 4380 49532
rect 4436 49530 4460 49532
rect 4516 49530 4522 49532
rect 4276 49478 4278 49530
rect 4458 49478 4460 49530
rect 4214 49476 4220 49478
rect 4276 49476 4300 49478
rect 4356 49476 4380 49478
rect 4436 49476 4460 49478
rect 4516 49476 4522 49478
rect 4214 49456 4522 49476
rect 4214 48444 4522 48464
rect 4214 48442 4220 48444
rect 4276 48442 4300 48444
rect 4356 48442 4380 48444
rect 4436 48442 4460 48444
rect 4516 48442 4522 48444
rect 4276 48390 4278 48442
rect 4458 48390 4460 48442
rect 4214 48388 4220 48390
rect 4276 48388 4300 48390
rect 4356 48388 4380 48390
rect 4436 48388 4460 48390
rect 4516 48388 4522 48390
rect 4214 48368 4522 48388
rect 4214 47356 4522 47376
rect 4214 47354 4220 47356
rect 4276 47354 4300 47356
rect 4356 47354 4380 47356
rect 4436 47354 4460 47356
rect 4516 47354 4522 47356
rect 4276 47302 4278 47354
rect 4458 47302 4460 47354
rect 4214 47300 4220 47302
rect 4276 47300 4300 47302
rect 4356 47300 4380 47302
rect 4436 47300 4460 47302
rect 4516 47300 4522 47302
rect 4214 47280 4522 47300
rect 4214 46268 4522 46288
rect 4214 46266 4220 46268
rect 4276 46266 4300 46268
rect 4356 46266 4380 46268
rect 4436 46266 4460 46268
rect 4516 46266 4522 46268
rect 4276 46214 4278 46266
rect 4458 46214 4460 46266
rect 4214 46212 4220 46214
rect 4276 46212 4300 46214
rect 4356 46212 4380 46214
rect 4436 46212 4460 46214
rect 4516 46212 4522 46214
rect 4214 46192 4522 46212
rect 4214 45180 4522 45200
rect 4214 45178 4220 45180
rect 4276 45178 4300 45180
rect 4356 45178 4380 45180
rect 4436 45178 4460 45180
rect 4516 45178 4522 45180
rect 4276 45126 4278 45178
rect 4458 45126 4460 45178
rect 4214 45124 4220 45126
rect 4276 45124 4300 45126
rect 4356 45124 4380 45126
rect 4436 45124 4460 45126
rect 4516 45124 4522 45126
rect 4214 45104 4522 45124
rect 4214 44092 4522 44112
rect 4214 44090 4220 44092
rect 4276 44090 4300 44092
rect 4356 44090 4380 44092
rect 4436 44090 4460 44092
rect 4516 44090 4522 44092
rect 4276 44038 4278 44090
rect 4458 44038 4460 44090
rect 4214 44036 4220 44038
rect 4276 44036 4300 44038
rect 4356 44036 4380 44038
rect 4436 44036 4460 44038
rect 4516 44036 4522 44038
rect 4214 44016 4522 44036
rect 4214 43004 4522 43024
rect 4214 43002 4220 43004
rect 4276 43002 4300 43004
rect 4356 43002 4380 43004
rect 4436 43002 4460 43004
rect 4516 43002 4522 43004
rect 4276 42950 4278 43002
rect 4458 42950 4460 43002
rect 4214 42948 4220 42950
rect 4276 42948 4300 42950
rect 4356 42948 4380 42950
rect 4436 42948 4460 42950
rect 4516 42948 4522 42950
rect 4214 42928 4522 42948
rect 4214 41916 4522 41936
rect 4214 41914 4220 41916
rect 4276 41914 4300 41916
rect 4356 41914 4380 41916
rect 4436 41914 4460 41916
rect 4516 41914 4522 41916
rect 4276 41862 4278 41914
rect 4458 41862 4460 41914
rect 4214 41860 4220 41862
rect 4276 41860 4300 41862
rect 4356 41860 4380 41862
rect 4436 41860 4460 41862
rect 4516 41860 4522 41862
rect 4214 41840 4522 41860
rect 4214 40828 4522 40848
rect 4214 40826 4220 40828
rect 4276 40826 4300 40828
rect 4356 40826 4380 40828
rect 4436 40826 4460 40828
rect 4516 40826 4522 40828
rect 4276 40774 4278 40826
rect 4458 40774 4460 40826
rect 4214 40772 4220 40774
rect 4276 40772 4300 40774
rect 4356 40772 4380 40774
rect 4436 40772 4460 40774
rect 4516 40772 4522 40774
rect 4214 40752 4522 40772
rect 4214 39740 4522 39760
rect 4214 39738 4220 39740
rect 4276 39738 4300 39740
rect 4356 39738 4380 39740
rect 4436 39738 4460 39740
rect 4516 39738 4522 39740
rect 4276 39686 4278 39738
rect 4458 39686 4460 39738
rect 4214 39684 4220 39686
rect 4276 39684 4300 39686
rect 4356 39684 4380 39686
rect 4436 39684 4460 39686
rect 4516 39684 4522 39686
rect 4214 39664 4522 39684
rect 4214 38652 4522 38672
rect 4214 38650 4220 38652
rect 4276 38650 4300 38652
rect 4356 38650 4380 38652
rect 4436 38650 4460 38652
rect 4516 38650 4522 38652
rect 4276 38598 4278 38650
rect 4458 38598 4460 38650
rect 4214 38596 4220 38598
rect 4276 38596 4300 38598
rect 4356 38596 4380 38598
rect 4436 38596 4460 38598
rect 4516 38596 4522 38598
rect 4214 38576 4522 38596
rect 4214 37564 4522 37584
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37488 4522 37508
rect 4214 36476 4522 36496
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36400 4522 36420
rect 4214 35388 4522 35408
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35312 4522 35332
rect 4214 34300 4522 34320
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34224 4522 34244
rect 4214 33212 4522 33232
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33136 4522 33156
rect 4214 32124 4522 32144
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32048 4522 32068
rect 4214 31036 4522 31056
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30960 4522 30980
rect 4214 29948 4522 29968
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29872 4522 29892
rect 4214 28860 4522 28880
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28784 4522 28804
rect 4214 27772 4522 27792
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27696 4522 27716
rect 4214 26684 4522 26704
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26608 4522 26628
rect 4214 25596 4522 25616
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25520 4522 25540
rect 4214 24508 4522 24528
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24432 4522 24452
rect 4214 23420 4522 23440
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23344 4522 23364
rect 4214 22332 4522 22352
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22256 4522 22276
rect 4214 21244 4522 21264
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21168 4522 21188
rect 4214 20156 4522 20176
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20080 4522 20100
rect 4214 19068 4522 19088
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 18992 4522 19012
rect 4214 17980 4522 18000
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17904 4522 17924
rect 4214 16892 4522 16912
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16816 4522 16836
rect 4214 15804 4522 15824
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15728 4522 15748
rect 4214 14716 4522 14736
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14640 4522 14660
rect 4214 13628 4522 13648
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13552 4522 13572
rect 4214 12540 4522 12560
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12464 4522 12484
rect 3056 11824 3108 11830
rect 3056 11766 3108 11772
rect 4214 11452 4522 11472
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11376 4522 11396
rect 4214 10364 4522 10384
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10288 4522 10308
rect 4214 9276 4522 9296
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9200 4522 9220
rect 4214 8188 4522 8208
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8112 4522 8132
rect 4214 7100 4522 7120
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7024 4522 7044
rect 4214 6012 4522 6032
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5936 4522 5956
rect 4214 4924 4522 4944
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4848 4522 4868
rect 4214 3836 4522 3856
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3760 4522 3780
rect 4214 2748 4522 2768
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2672 4522 2692
rect 4632 2514 4660 59706
rect 19574 58780 19882 58800
rect 19574 58778 19580 58780
rect 19636 58778 19660 58780
rect 19716 58778 19740 58780
rect 19796 58778 19820 58780
rect 19876 58778 19882 58780
rect 19636 58726 19638 58778
rect 19818 58726 19820 58778
rect 19574 58724 19580 58726
rect 19636 58724 19660 58726
rect 19716 58724 19740 58726
rect 19796 58724 19820 58726
rect 19876 58724 19882 58726
rect 19574 58704 19882 58724
rect 19574 57692 19882 57712
rect 19574 57690 19580 57692
rect 19636 57690 19660 57692
rect 19716 57690 19740 57692
rect 19796 57690 19820 57692
rect 19876 57690 19882 57692
rect 19636 57638 19638 57690
rect 19818 57638 19820 57690
rect 19574 57636 19580 57638
rect 19636 57636 19660 57638
rect 19716 57636 19740 57638
rect 19796 57636 19820 57638
rect 19876 57636 19882 57638
rect 19574 57616 19882 57636
rect 19574 56604 19882 56624
rect 19574 56602 19580 56604
rect 19636 56602 19660 56604
rect 19716 56602 19740 56604
rect 19796 56602 19820 56604
rect 19876 56602 19882 56604
rect 19636 56550 19638 56602
rect 19818 56550 19820 56602
rect 19574 56548 19580 56550
rect 19636 56548 19660 56550
rect 19716 56548 19740 56550
rect 19796 56548 19820 56550
rect 19876 56548 19882 56550
rect 19574 56528 19882 56548
rect 19574 55516 19882 55536
rect 19574 55514 19580 55516
rect 19636 55514 19660 55516
rect 19716 55514 19740 55516
rect 19796 55514 19820 55516
rect 19876 55514 19882 55516
rect 19636 55462 19638 55514
rect 19818 55462 19820 55514
rect 19574 55460 19580 55462
rect 19636 55460 19660 55462
rect 19716 55460 19740 55462
rect 19796 55460 19820 55462
rect 19876 55460 19882 55462
rect 19574 55440 19882 55460
rect 19574 54428 19882 54448
rect 19574 54426 19580 54428
rect 19636 54426 19660 54428
rect 19716 54426 19740 54428
rect 19796 54426 19820 54428
rect 19876 54426 19882 54428
rect 19636 54374 19638 54426
rect 19818 54374 19820 54426
rect 19574 54372 19580 54374
rect 19636 54372 19660 54374
rect 19716 54372 19740 54374
rect 19796 54372 19820 54374
rect 19876 54372 19882 54374
rect 19574 54352 19882 54372
rect 19574 53340 19882 53360
rect 19574 53338 19580 53340
rect 19636 53338 19660 53340
rect 19716 53338 19740 53340
rect 19796 53338 19820 53340
rect 19876 53338 19882 53340
rect 19636 53286 19638 53338
rect 19818 53286 19820 53338
rect 19574 53284 19580 53286
rect 19636 53284 19660 53286
rect 19716 53284 19740 53286
rect 19796 53284 19820 53286
rect 19876 53284 19882 53286
rect 19574 53264 19882 53284
rect 19574 52252 19882 52272
rect 19574 52250 19580 52252
rect 19636 52250 19660 52252
rect 19716 52250 19740 52252
rect 19796 52250 19820 52252
rect 19876 52250 19882 52252
rect 19636 52198 19638 52250
rect 19818 52198 19820 52250
rect 19574 52196 19580 52198
rect 19636 52196 19660 52198
rect 19716 52196 19740 52198
rect 19796 52196 19820 52198
rect 19876 52196 19882 52198
rect 19574 52176 19882 52196
rect 19574 51164 19882 51184
rect 19574 51162 19580 51164
rect 19636 51162 19660 51164
rect 19716 51162 19740 51164
rect 19796 51162 19820 51164
rect 19876 51162 19882 51164
rect 19636 51110 19638 51162
rect 19818 51110 19820 51162
rect 19574 51108 19580 51110
rect 19636 51108 19660 51110
rect 19716 51108 19740 51110
rect 19796 51108 19820 51110
rect 19876 51108 19882 51110
rect 19574 51088 19882 51108
rect 19574 50076 19882 50096
rect 19574 50074 19580 50076
rect 19636 50074 19660 50076
rect 19716 50074 19740 50076
rect 19796 50074 19820 50076
rect 19876 50074 19882 50076
rect 19636 50022 19638 50074
rect 19818 50022 19820 50074
rect 19574 50020 19580 50022
rect 19636 50020 19660 50022
rect 19716 50020 19740 50022
rect 19796 50020 19820 50022
rect 19876 50020 19882 50022
rect 19574 50000 19882 50020
rect 19574 48988 19882 49008
rect 19574 48986 19580 48988
rect 19636 48986 19660 48988
rect 19716 48986 19740 48988
rect 19796 48986 19820 48988
rect 19876 48986 19882 48988
rect 19636 48934 19638 48986
rect 19818 48934 19820 48986
rect 19574 48932 19580 48934
rect 19636 48932 19660 48934
rect 19716 48932 19740 48934
rect 19796 48932 19820 48934
rect 19876 48932 19882 48934
rect 19574 48912 19882 48932
rect 19574 47900 19882 47920
rect 19574 47898 19580 47900
rect 19636 47898 19660 47900
rect 19716 47898 19740 47900
rect 19796 47898 19820 47900
rect 19876 47898 19882 47900
rect 19636 47846 19638 47898
rect 19818 47846 19820 47898
rect 19574 47844 19580 47846
rect 19636 47844 19660 47846
rect 19716 47844 19740 47846
rect 19796 47844 19820 47846
rect 19876 47844 19882 47846
rect 19574 47824 19882 47844
rect 19574 46812 19882 46832
rect 19574 46810 19580 46812
rect 19636 46810 19660 46812
rect 19716 46810 19740 46812
rect 19796 46810 19820 46812
rect 19876 46810 19882 46812
rect 19636 46758 19638 46810
rect 19818 46758 19820 46810
rect 19574 46756 19580 46758
rect 19636 46756 19660 46758
rect 19716 46756 19740 46758
rect 19796 46756 19820 46758
rect 19876 46756 19882 46758
rect 19574 46736 19882 46756
rect 19574 45724 19882 45744
rect 19574 45722 19580 45724
rect 19636 45722 19660 45724
rect 19716 45722 19740 45724
rect 19796 45722 19820 45724
rect 19876 45722 19882 45724
rect 19636 45670 19638 45722
rect 19818 45670 19820 45722
rect 19574 45668 19580 45670
rect 19636 45668 19660 45670
rect 19716 45668 19740 45670
rect 19796 45668 19820 45670
rect 19876 45668 19882 45670
rect 19574 45648 19882 45668
rect 19574 44636 19882 44656
rect 19574 44634 19580 44636
rect 19636 44634 19660 44636
rect 19716 44634 19740 44636
rect 19796 44634 19820 44636
rect 19876 44634 19882 44636
rect 19636 44582 19638 44634
rect 19818 44582 19820 44634
rect 19574 44580 19580 44582
rect 19636 44580 19660 44582
rect 19716 44580 19740 44582
rect 19796 44580 19820 44582
rect 19876 44580 19882 44582
rect 19574 44560 19882 44580
rect 19574 43548 19882 43568
rect 19574 43546 19580 43548
rect 19636 43546 19660 43548
rect 19716 43546 19740 43548
rect 19796 43546 19820 43548
rect 19876 43546 19882 43548
rect 19636 43494 19638 43546
rect 19818 43494 19820 43546
rect 19574 43492 19580 43494
rect 19636 43492 19660 43494
rect 19716 43492 19740 43494
rect 19796 43492 19820 43494
rect 19876 43492 19882 43494
rect 19574 43472 19882 43492
rect 19574 42460 19882 42480
rect 19574 42458 19580 42460
rect 19636 42458 19660 42460
rect 19716 42458 19740 42460
rect 19796 42458 19820 42460
rect 19876 42458 19882 42460
rect 19636 42406 19638 42458
rect 19818 42406 19820 42458
rect 19574 42404 19580 42406
rect 19636 42404 19660 42406
rect 19716 42404 19740 42406
rect 19796 42404 19820 42406
rect 19876 42404 19882 42406
rect 19574 42384 19882 42404
rect 19574 41372 19882 41392
rect 19574 41370 19580 41372
rect 19636 41370 19660 41372
rect 19716 41370 19740 41372
rect 19796 41370 19820 41372
rect 19876 41370 19882 41372
rect 19636 41318 19638 41370
rect 19818 41318 19820 41370
rect 19574 41316 19580 41318
rect 19636 41316 19660 41318
rect 19716 41316 19740 41318
rect 19796 41316 19820 41318
rect 19876 41316 19882 41318
rect 19574 41296 19882 41316
rect 19574 40284 19882 40304
rect 19574 40282 19580 40284
rect 19636 40282 19660 40284
rect 19716 40282 19740 40284
rect 19796 40282 19820 40284
rect 19876 40282 19882 40284
rect 19636 40230 19638 40282
rect 19818 40230 19820 40282
rect 19574 40228 19580 40230
rect 19636 40228 19660 40230
rect 19716 40228 19740 40230
rect 19796 40228 19820 40230
rect 19876 40228 19882 40230
rect 19574 40208 19882 40228
rect 19574 39196 19882 39216
rect 19574 39194 19580 39196
rect 19636 39194 19660 39196
rect 19716 39194 19740 39196
rect 19796 39194 19820 39196
rect 19876 39194 19882 39196
rect 19636 39142 19638 39194
rect 19818 39142 19820 39194
rect 19574 39140 19580 39142
rect 19636 39140 19660 39142
rect 19716 39140 19740 39142
rect 19796 39140 19820 39142
rect 19876 39140 19882 39142
rect 19574 39120 19882 39140
rect 19574 38108 19882 38128
rect 19574 38106 19580 38108
rect 19636 38106 19660 38108
rect 19716 38106 19740 38108
rect 19796 38106 19820 38108
rect 19876 38106 19882 38108
rect 19636 38054 19638 38106
rect 19818 38054 19820 38106
rect 19574 38052 19580 38054
rect 19636 38052 19660 38054
rect 19716 38052 19740 38054
rect 19796 38052 19820 38054
rect 19876 38052 19882 38054
rect 19574 38032 19882 38052
rect 19574 37020 19882 37040
rect 19574 37018 19580 37020
rect 19636 37018 19660 37020
rect 19716 37018 19740 37020
rect 19796 37018 19820 37020
rect 19876 37018 19882 37020
rect 19636 36966 19638 37018
rect 19818 36966 19820 37018
rect 19574 36964 19580 36966
rect 19636 36964 19660 36966
rect 19716 36964 19740 36966
rect 19796 36964 19820 36966
rect 19876 36964 19882 36966
rect 19574 36944 19882 36964
rect 19574 35932 19882 35952
rect 19574 35930 19580 35932
rect 19636 35930 19660 35932
rect 19716 35930 19740 35932
rect 19796 35930 19820 35932
rect 19876 35930 19882 35932
rect 19636 35878 19638 35930
rect 19818 35878 19820 35930
rect 19574 35876 19580 35878
rect 19636 35876 19660 35878
rect 19716 35876 19740 35878
rect 19796 35876 19820 35878
rect 19876 35876 19882 35878
rect 19574 35856 19882 35876
rect 19574 34844 19882 34864
rect 19574 34842 19580 34844
rect 19636 34842 19660 34844
rect 19716 34842 19740 34844
rect 19796 34842 19820 34844
rect 19876 34842 19882 34844
rect 19636 34790 19638 34842
rect 19818 34790 19820 34842
rect 19574 34788 19580 34790
rect 19636 34788 19660 34790
rect 19716 34788 19740 34790
rect 19796 34788 19820 34790
rect 19876 34788 19882 34790
rect 19574 34768 19882 34788
rect 19574 33756 19882 33776
rect 19574 33754 19580 33756
rect 19636 33754 19660 33756
rect 19716 33754 19740 33756
rect 19796 33754 19820 33756
rect 19876 33754 19882 33756
rect 19636 33702 19638 33754
rect 19818 33702 19820 33754
rect 19574 33700 19580 33702
rect 19636 33700 19660 33702
rect 19716 33700 19740 33702
rect 19796 33700 19820 33702
rect 19876 33700 19882 33702
rect 19574 33680 19882 33700
rect 19574 32668 19882 32688
rect 19574 32666 19580 32668
rect 19636 32666 19660 32668
rect 19716 32666 19740 32668
rect 19796 32666 19820 32668
rect 19876 32666 19882 32668
rect 19636 32614 19638 32666
rect 19818 32614 19820 32666
rect 19574 32612 19580 32614
rect 19636 32612 19660 32614
rect 19716 32612 19740 32614
rect 19796 32612 19820 32614
rect 19876 32612 19882 32614
rect 19574 32592 19882 32612
rect 19574 31580 19882 31600
rect 19574 31578 19580 31580
rect 19636 31578 19660 31580
rect 19716 31578 19740 31580
rect 19796 31578 19820 31580
rect 19876 31578 19882 31580
rect 19636 31526 19638 31578
rect 19818 31526 19820 31578
rect 19574 31524 19580 31526
rect 19636 31524 19660 31526
rect 19716 31524 19740 31526
rect 19796 31524 19820 31526
rect 19876 31524 19882 31526
rect 19574 31504 19882 31524
rect 19574 30492 19882 30512
rect 19574 30490 19580 30492
rect 19636 30490 19660 30492
rect 19716 30490 19740 30492
rect 19796 30490 19820 30492
rect 19876 30490 19882 30492
rect 19636 30438 19638 30490
rect 19818 30438 19820 30490
rect 19574 30436 19580 30438
rect 19636 30436 19660 30438
rect 19716 30436 19740 30438
rect 19796 30436 19820 30438
rect 19876 30436 19882 30438
rect 19574 30416 19882 30436
rect 19574 29404 19882 29424
rect 19574 29402 19580 29404
rect 19636 29402 19660 29404
rect 19716 29402 19740 29404
rect 19796 29402 19820 29404
rect 19876 29402 19882 29404
rect 19636 29350 19638 29402
rect 19818 29350 19820 29402
rect 19574 29348 19580 29350
rect 19636 29348 19660 29350
rect 19716 29348 19740 29350
rect 19796 29348 19820 29350
rect 19876 29348 19882 29350
rect 19574 29328 19882 29348
rect 19574 28316 19882 28336
rect 19574 28314 19580 28316
rect 19636 28314 19660 28316
rect 19716 28314 19740 28316
rect 19796 28314 19820 28316
rect 19876 28314 19882 28316
rect 19636 28262 19638 28314
rect 19818 28262 19820 28314
rect 19574 28260 19580 28262
rect 19636 28260 19660 28262
rect 19716 28260 19740 28262
rect 19796 28260 19820 28262
rect 19876 28260 19882 28262
rect 19574 28240 19882 28260
rect 19574 27228 19882 27248
rect 19574 27226 19580 27228
rect 19636 27226 19660 27228
rect 19716 27226 19740 27228
rect 19796 27226 19820 27228
rect 19876 27226 19882 27228
rect 19636 27174 19638 27226
rect 19818 27174 19820 27226
rect 19574 27172 19580 27174
rect 19636 27172 19660 27174
rect 19716 27172 19740 27174
rect 19796 27172 19820 27174
rect 19876 27172 19882 27174
rect 19574 27152 19882 27172
rect 19574 26140 19882 26160
rect 19574 26138 19580 26140
rect 19636 26138 19660 26140
rect 19716 26138 19740 26140
rect 19796 26138 19820 26140
rect 19876 26138 19882 26140
rect 19636 26086 19638 26138
rect 19818 26086 19820 26138
rect 19574 26084 19580 26086
rect 19636 26084 19660 26086
rect 19716 26084 19740 26086
rect 19796 26084 19820 26086
rect 19876 26084 19882 26086
rect 19574 26064 19882 26084
rect 19574 25052 19882 25072
rect 19574 25050 19580 25052
rect 19636 25050 19660 25052
rect 19716 25050 19740 25052
rect 19796 25050 19820 25052
rect 19876 25050 19882 25052
rect 19636 24998 19638 25050
rect 19818 24998 19820 25050
rect 19574 24996 19580 24998
rect 19636 24996 19660 24998
rect 19716 24996 19740 24998
rect 19796 24996 19820 24998
rect 19876 24996 19882 24998
rect 19574 24976 19882 24996
rect 19574 23964 19882 23984
rect 19574 23962 19580 23964
rect 19636 23962 19660 23964
rect 19716 23962 19740 23964
rect 19796 23962 19820 23964
rect 19876 23962 19882 23964
rect 19636 23910 19638 23962
rect 19818 23910 19820 23962
rect 19574 23908 19580 23910
rect 19636 23908 19660 23910
rect 19716 23908 19740 23910
rect 19796 23908 19820 23910
rect 19876 23908 19882 23910
rect 19574 23888 19882 23908
rect 19574 22876 19882 22896
rect 19574 22874 19580 22876
rect 19636 22874 19660 22876
rect 19716 22874 19740 22876
rect 19796 22874 19820 22876
rect 19876 22874 19882 22876
rect 19636 22822 19638 22874
rect 19818 22822 19820 22874
rect 19574 22820 19580 22822
rect 19636 22820 19660 22822
rect 19716 22820 19740 22822
rect 19796 22820 19820 22822
rect 19876 22820 19882 22822
rect 19574 22800 19882 22820
rect 19574 21788 19882 21808
rect 19574 21786 19580 21788
rect 19636 21786 19660 21788
rect 19716 21786 19740 21788
rect 19796 21786 19820 21788
rect 19876 21786 19882 21788
rect 19636 21734 19638 21786
rect 19818 21734 19820 21786
rect 19574 21732 19580 21734
rect 19636 21732 19660 21734
rect 19716 21732 19740 21734
rect 19796 21732 19820 21734
rect 19876 21732 19882 21734
rect 19574 21712 19882 21732
rect 19574 20700 19882 20720
rect 19574 20698 19580 20700
rect 19636 20698 19660 20700
rect 19716 20698 19740 20700
rect 19796 20698 19820 20700
rect 19876 20698 19882 20700
rect 19636 20646 19638 20698
rect 19818 20646 19820 20698
rect 19574 20644 19580 20646
rect 19636 20644 19660 20646
rect 19716 20644 19740 20646
rect 19796 20644 19820 20646
rect 19876 20644 19882 20646
rect 19574 20624 19882 20644
rect 19574 19612 19882 19632
rect 19574 19610 19580 19612
rect 19636 19610 19660 19612
rect 19716 19610 19740 19612
rect 19796 19610 19820 19612
rect 19876 19610 19882 19612
rect 19636 19558 19638 19610
rect 19818 19558 19820 19610
rect 19574 19556 19580 19558
rect 19636 19556 19660 19558
rect 19716 19556 19740 19558
rect 19796 19556 19820 19558
rect 19876 19556 19882 19558
rect 19574 19536 19882 19556
rect 19574 18524 19882 18544
rect 19574 18522 19580 18524
rect 19636 18522 19660 18524
rect 19716 18522 19740 18524
rect 19796 18522 19820 18524
rect 19876 18522 19882 18524
rect 19636 18470 19638 18522
rect 19818 18470 19820 18522
rect 19574 18468 19580 18470
rect 19636 18468 19660 18470
rect 19716 18468 19740 18470
rect 19796 18468 19820 18470
rect 19876 18468 19882 18470
rect 19574 18448 19882 18468
rect 19574 17436 19882 17456
rect 19574 17434 19580 17436
rect 19636 17434 19660 17436
rect 19716 17434 19740 17436
rect 19796 17434 19820 17436
rect 19876 17434 19882 17436
rect 19636 17382 19638 17434
rect 19818 17382 19820 17434
rect 19574 17380 19580 17382
rect 19636 17380 19660 17382
rect 19716 17380 19740 17382
rect 19796 17380 19820 17382
rect 19876 17380 19882 17382
rect 19574 17360 19882 17380
rect 19574 16348 19882 16368
rect 19574 16346 19580 16348
rect 19636 16346 19660 16348
rect 19716 16346 19740 16348
rect 19796 16346 19820 16348
rect 19876 16346 19882 16348
rect 19636 16294 19638 16346
rect 19818 16294 19820 16346
rect 19574 16292 19580 16294
rect 19636 16292 19660 16294
rect 19716 16292 19740 16294
rect 19796 16292 19820 16294
rect 19876 16292 19882 16294
rect 19574 16272 19882 16292
rect 19574 15260 19882 15280
rect 19574 15258 19580 15260
rect 19636 15258 19660 15260
rect 19716 15258 19740 15260
rect 19796 15258 19820 15260
rect 19876 15258 19882 15260
rect 19636 15206 19638 15258
rect 19818 15206 19820 15258
rect 19574 15204 19580 15206
rect 19636 15204 19660 15206
rect 19716 15204 19740 15206
rect 19796 15204 19820 15206
rect 19876 15204 19882 15206
rect 19574 15184 19882 15204
rect 19574 14172 19882 14192
rect 19574 14170 19580 14172
rect 19636 14170 19660 14172
rect 19716 14170 19740 14172
rect 19796 14170 19820 14172
rect 19876 14170 19882 14172
rect 19636 14118 19638 14170
rect 19818 14118 19820 14170
rect 19574 14116 19580 14118
rect 19636 14116 19660 14118
rect 19716 14116 19740 14118
rect 19796 14116 19820 14118
rect 19876 14116 19882 14118
rect 19574 14096 19882 14116
rect 19574 13084 19882 13104
rect 19574 13082 19580 13084
rect 19636 13082 19660 13084
rect 19716 13082 19740 13084
rect 19796 13082 19820 13084
rect 19876 13082 19882 13084
rect 19636 13030 19638 13082
rect 19818 13030 19820 13082
rect 19574 13028 19580 13030
rect 19636 13028 19660 13030
rect 19716 13028 19740 13030
rect 19796 13028 19820 13030
rect 19876 13028 19882 13030
rect 19574 13008 19882 13028
rect 18328 12164 18380 12170
rect 18328 12106 18380 12112
rect 12440 3528 12492 3534
rect 12440 3470 12492 3476
rect 11520 3188 11572 3194
rect 11520 3130 11572 3136
rect 4620 2508 4672 2514
rect 4620 2450 4672 2456
rect 11532 2446 11560 3130
rect 12452 2582 12480 3470
rect 16212 3392 16264 3398
rect 16212 3334 16264 3340
rect 12440 2576 12492 2582
rect 12440 2518 12492 2524
rect 16224 2446 16252 3334
rect 18340 2650 18368 12106
rect 19574 11996 19882 12016
rect 19574 11994 19580 11996
rect 19636 11994 19660 11996
rect 19716 11994 19740 11996
rect 19796 11994 19820 11996
rect 19876 11994 19882 11996
rect 19636 11942 19638 11994
rect 19818 11942 19820 11994
rect 19574 11940 19580 11942
rect 19636 11940 19660 11942
rect 19716 11940 19740 11942
rect 19796 11940 19820 11942
rect 19876 11940 19882 11942
rect 19574 11920 19882 11940
rect 19574 10908 19882 10928
rect 19574 10906 19580 10908
rect 19636 10906 19660 10908
rect 19716 10906 19740 10908
rect 19796 10906 19820 10908
rect 19876 10906 19882 10908
rect 19636 10854 19638 10906
rect 19818 10854 19820 10906
rect 19574 10852 19580 10854
rect 19636 10852 19660 10854
rect 19716 10852 19740 10854
rect 19796 10852 19820 10854
rect 19876 10852 19882 10854
rect 19574 10832 19882 10852
rect 19574 9820 19882 9840
rect 19574 9818 19580 9820
rect 19636 9818 19660 9820
rect 19716 9818 19740 9820
rect 19796 9818 19820 9820
rect 19876 9818 19882 9820
rect 19636 9766 19638 9818
rect 19818 9766 19820 9818
rect 19574 9764 19580 9766
rect 19636 9764 19660 9766
rect 19716 9764 19740 9766
rect 19796 9764 19820 9766
rect 19876 9764 19882 9766
rect 19574 9744 19882 9764
rect 19574 8732 19882 8752
rect 19574 8730 19580 8732
rect 19636 8730 19660 8732
rect 19716 8730 19740 8732
rect 19796 8730 19820 8732
rect 19876 8730 19882 8732
rect 19636 8678 19638 8730
rect 19818 8678 19820 8730
rect 19574 8676 19580 8678
rect 19636 8676 19660 8678
rect 19716 8676 19740 8678
rect 19796 8676 19820 8678
rect 19876 8676 19882 8678
rect 19574 8656 19882 8676
rect 19574 7644 19882 7664
rect 19574 7642 19580 7644
rect 19636 7642 19660 7644
rect 19716 7642 19740 7644
rect 19796 7642 19820 7644
rect 19876 7642 19882 7644
rect 19636 7590 19638 7642
rect 19818 7590 19820 7642
rect 19574 7588 19580 7590
rect 19636 7588 19660 7590
rect 19716 7588 19740 7590
rect 19796 7588 19820 7590
rect 19876 7588 19882 7590
rect 19574 7568 19882 7588
rect 19574 6556 19882 6576
rect 19574 6554 19580 6556
rect 19636 6554 19660 6556
rect 19716 6554 19740 6556
rect 19796 6554 19820 6556
rect 19876 6554 19882 6556
rect 19636 6502 19638 6554
rect 19818 6502 19820 6554
rect 19574 6500 19580 6502
rect 19636 6500 19660 6502
rect 19716 6500 19740 6502
rect 19796 6500 19820 6502
rect 19876 6500 19882 6502
rect 19574 6480 19882 6500
rect 19574 5468 19882 5488
rect 19574 5466 19580 5468
rect 19636 5466 19660 5468
rect 19716 5466 19740 5468
rect 19796 5466 19820 5468
rect 19876 5466 19882 5468
rect 19636 5414 19638 5466
rect 19818 5414 19820 5466
rect 19574 5412 19580 5414
rect 19636 5412 19660 5414
rect 19716 5412 19740 5414
rect 19796 5412 19820 5414
rect 19876 5412 19882 5414
rect 19574 5392 19882 5412
rect 19574 4380 19882 4400
rect 19574 4378 19580 4380
rect 19636 4378 19660 4380
rect 19716 4378 19740 4380
rect 19796 4378 19820 4380
rect 19876 4378 19882 4380
rect 19636 4326 19638 4378
rect 19818 4326 19820 4378
rect 19574 4324 19580 4326
rect 19636 4324 19660 4326
rect 19716 4324 19740 4326
rect 19796 4324 19820 4326
rect 19876 4324 19882 4326
rect 19574 4304 19882 4324
rect 19574 3292 19882 3312
rect 19574 3290 19580 3292
rect 19636 3290 19660 3292
rect 19716 3290 19740 3292
rect 19796 3290 19820 3292
rect 19876 3290 19882 3292
rect 19636 3238 19638 3290
rect 19818 3238 19820 3290
rect 19574 3236 19580 3238
rect 19636 3236 19660 3238
rect 19716 3236 19740 3238
rect 19796 3236 19820 3238
rect 19876 3236 19882 3238
rect 19574 3216 19882 3236
rect 18328 2644 18380 2650
rect 18328 2586 18380 2592
rect 19996 2514 20024 59978
rect 35348 59968 35400 59974
rect 35348 59910 35400 59916
rect 33140 59764 33192 59770
rect 33140 59706 33192 59712
rect 29920 7404 29972 7410
rect 29920 7346 29972 7352
rect 29932 2650 29960 7346
rect 33152 2650 33180 59706
rect 34934 59324 35242 59344
rect 34934 59322 34940 59324
rect 34996 59322 35020 59324
rect 35076 59322 35100 59324
rect 35156 59322 35180 59324
rect 35236 59322 35242 59324
rect 34996 59270 34998 59322
rect 35178 59270 35180 59322
rect 34934 59268 34940 59270
rect 34996 59268 35020 59270
rect 35076 59268 35100 59270
rect 35156 59268 35180 59270
rect 35236 59268 35242 59270
rect 34934 59248 35242 59268
rect 34934 58236 35242 58256
rect 34934 58234 34940 58236
rect 34996 58234 35020 58236
rect 35076 58234 35100 58236
rect 35156 58234 35180 58236
rect 35236 58234 35242 58236
rect 34996 58182 34998 58234
rect 35178 58182 35180 58234
rect 34934 58180 34940 58182
rect 34996 58180 35020 58182
rect 35076 58180 35100 58182
rect 35156 58180 35180 58182
rect 35236 58180 35242 58182
rect 34934 58160 35242 58180
rect 34934 57148 35242 57168
rect 34934 57146 34940 57148
rect 34996 57146 35020 57148
rect 35076 57146 35100 57148
rect 35156 57146 35180 57148
rect 35236 57146 35242 57148
rect 34996 57094 34998 57146
rect 35178 57094 35180 57146
rect 34934 57092 34940 57094
rect 34996 57092 35020 57094
rect 35076 57092 35100 57094
rect 35156 57092 35180 57094
rect 35236 57092 35242 57094
rect 34934 57072 35242 57092
rect 34934 56060 35242 56080
rect 34934 56058 34940 56060
rect 34996 56058 35020 56060
rect 35076 56058 35100 56060
rect 35156 56058 35180 56060
rect 35236 56058 35242 56060
rect 34996 56006 34998 56058
rect 35178 56006 35180 56058
rect 34934 56004 34940 56006
rect 34996 56004 35020 56006
rect 35076 56004 35100 56006
rect 35156 56004 35180 56006
rect 35236 56004 35242 56006
rect 34934 55984 35242 56004
rect 34934 54972 35242 54992
rect 34934 54970 34940 54972
rect 34996 54970 35020 54972
rect 35076 54970 35100 54972
rect 35156 54970 35180 54972
rect 35236 54970 35242 54972
rect 34996 54918 34998 54970
rect 35178 54918 35180 54970
rect 34934 54916 34940 54918
rect 34996 54916 35020 54918
rect 35076 54916 35100 54918
rect 35156 54916 35180 54918
rect 35236 54916 35242 54918
rect 34934 54896 35242 54916
rect 34934 53884 35242 53904
rect 34934 53882 34940 53884
rect 34996 53882 35020 53884
rect 35076 53882 35100 53884
rect 35156 53882 35180 53884
rect 35236 53882 35242 53884
rect 34996 53830 34998 53882
rect 35178 53830 35180 53882
rect 34934 53828 34940 53830
rect 34996 53828 35020 53830
rect 35076 53828 35100 53830
rect 35156 53828 35180 53830
rect 35236 53828 35242 53830
rect 34934 53808 35242 53828
rect 34934 52796 35242 52816
rect 34934 52794 34940 52796
rect 34996 52794 35020 52796
rect 35076 52794 35100 52796
rect 35156 52794 35180 52796
rect 35236 52794 35242 52796
rect 34996 52742 34998 52794
rect 35178 52742 35180 52794
rect 34934 52740 34940 52742
rect 34996 52740 35020 52742
rect 35076 52740 35100 52742
rect 35156 52740 35180 52742
rect 35236 52740 35242 52742
rect 34934 52720 35242 52740
rect 34934 51708 35242 51728
rect 34934 51706 34940 51708
rect 34996 51706 35020 51708
rect 35076 51706 35100 51708
rect 35156 51706 35180 51708
rect 35236 51706 35242 51708
rect 34996 51654 34998 51706
rect 35178 51654 35180 51706
rect 34934 51652 34940 51654
rect 34996 51652 35020 51654
rect 35076 51652 35100 51654
rect 35156 51652 35180 51654
rect 35236 51652 35242 51654
rect 34934 51632 35242 51652
rect 34934 50620 35242 50640
rect 34934 50618 34940 50620
rect 34996 50618 35020 50620
rect 35076 50618 35100 50620
rect 35156 50618 35180 50620
rect 35236 50618 35242 50620
rect 34996 50566 34998 50618
rect 35178 50566 35180 50618
rect 34934 50564 34940 50566
rect 34996 50564 35020 50566
rect 35076 50564 35100 50566
rect 35156 50564 35180 50566
rect 35236 50564 35242 50566
rect 34934 50544 35242 50564
rect 34934 49532 35242 49552
rect 34934 49530 34940 49532
rect 34996 49530 35020 49532
rect 35076 49530 35100 49532
rect 35156 49530 35180 49532
rect 35236 49530 35242 49532
rect 34996 49478 34998 49530
rect 35178 49478 35180 49530
rect 34934 49476 34940 49478
rect 34996 49476 35020 49478
rect 35076 49476 35100 49478
rect 35156 49476 35180 49478
rect 35236 49476 35242 49478
rect 34934 49456 35242 49476
rect 34934 48444 35242 48464
rect 34934 48442 34940 48444
rect 34996 48442 35020 48444
rect 35076 48442 35100 48444
rect 35156 48442 35180 48444
rect 35236 48442 35242 48444
rect 34996 48390 34998 48442
rect 35178 48390 35180 48442
rect 34934 48388 34940 48390
rect 34996 48388 35020 48390
rect 35076 48388 35100 48390
rect 35156 48388 35180 48390
rect 35236 48388 35242 48390
rect 34934 48368 35242 48388
rect 34934 47356 35242 47376
rect 34934 47354 34940 47356
rect 34996 47354 35020 47356
rect 35076 47354 35100 47356
rect 35156 47354 35180 47356
rect 35236 47354 35242 47356
rect 34996 47302 34998 47354
rect 35178 47302 35180 47354
rect 34934 47300 34940 47302
rect 34996 47300 35020 47302
rect 35076 47300 35100 47302
rect 35156 47300 35180 47302
rect 35236 47300 35242 47302
rect 34934 47280 35242 47300
rect 34934 46268 35242 46288
rect 34934 46266 34940 46268
rect 34996 46266 35020 46268
rect 35076 46266 35100 46268
rect 35156 46266 35180 46268
rect 35236 46266 35242 46268
rect 34996 46214 34998 46266
rect 35178 46214 35180 46266
rect 34934 46212 34940 46214
rect 34996 46212 35020 46214
rect 35076 46212 35100 46214
rect 35156 46212 35180 46214
rect 35236 46212 35242 46214
rect 34934 46192 35242 46212
rect 34934 45180 35242 45200
rect 34934 45178 34940 45180
rect 34996 45178 35020 45180
rect 35076 45178 35100 45180
rect 35156 45178 35180 45180
rect 35236 45178 35242 45180
rect 34996 45126 34998 45178
rect 35178 45126 35180 45178
rect 34934 45124 34940 45126
rect 34996 45124 35020 45126
rect 35076 45124 35100 45126
rect 35156 45124 35180 45126
rect 35236 45124 35242 45126
rect 34934 45104 35242 45124
rect 34934 44092 35242 44112
rect 34934 44090 34940 44092
rect 34996 44090 35020 44092
rect 35076 44090 35100 44092
rect 35156 44090 35180 44092
rect 35236 44090 35242 44092
rect 34996 44038 34998 44090
rect 35178 44038 35180 44090
rect 34934 44036 34940 44038
rect 34996 44036 35020 44038
rect 35076 44036 35100 44038
rect 35156 44036 35180 44038
rect 35236 44036 35242 44038
rect 34934 44016 35242 44036
rect 34934 43004 35242 43024
rect 34934 43002 34940 43004
rect 34996 43002 35020 43004
rect 35076 43002 35100 43004
rect 35156 43002 35180 43004
rect 35236 43002 35242 43004
rect 34996 42950 34998 43002
rect 35178 42950 35180 43002
rect 34934 42948 34940 42950
rect 34996 42948 35020 42950
rect 35076 42948 35100 42950
rect 35156 42948 35180 42950
rect 35236 42948 35242 42950
rect 34934 42928 35242 42948
rect 34934 41916 35242 41936
rect 34934 41914 34940 41916
rect 34996 41914 35020 41916
rect 35076 41914 35100 41916
rect 35156 41914 35180 41916
rect 35236 41914 35242 41916
rect 34996 41862 34998 41914
rect 35178 41862 35180 41914
rect 34934 41860 34940 41862
rect 34996 41860 35020 41862
rect 35076 41860 35100 41862
rect 35156 41860 35180 41862
rect 35236 41860 35242 41862
rect 34934 41840 35242 41860
rect 34934 40828 35242 40848
rect 34934 40826 34940 40828
rect 34996 40826 35020 40828
rect 35076 40826 35100 40828
rect 35156 40826 35180 40828
rect 35236 40826 35242 40828
rect 34996 40774 34998 40826
rect 35178 40774 35180 40826
rect 34934 40772 34940 40774
rect 34996 40772 35020 40774
rect 35076 40772 35100 40774
rect 35156 40772 35180 40774
rect 35236 40772 35242 40774
rect 34934 40752 35242 40772
rect 34934 39740 35242 39760
rect 34934 39738 34940 39740
rect 34996 39738 35020 39740
rect 35076 39738 35100 39740
rect 35156 39738 35180 39740
rect 35236 39738 35242 39740
rect 34996 39686 34998 39738
rect 35178 39686 35180 39738
rect 34934 39684 34940 39686
rect 34996 39684 35020 39686
rect 35076 39684 35100 39686
rect 35156 39684 35180 39686
rect 35236 39684 35242 39686
rect 34934 39664 35242 39684
rect 34934 38652 35242 38672
rect 34934 38650 34940 38652
rect 34996 38650 35020 38652
rect 35076 38650 35100 38652
rect 35156 38650 35180 38652
rect 35236 38650 35242 38652
rect 34996 38598 34998 38650
rect 35178 38598 35180 38650
rect 34934 38596 34940 38598
rect 34996 38596 35020 38598
rect 35076 38596 35100 38598
rect 35156 38596 35180 38598
rect 35236 38596 35242 38598
rect 34934 38576 35242 38596
rect 34934 37564 35242 37584
rect 34934 37562 34940 37564
rect 34996 37562 35020 37564
rect 35076 37562 35100 37564
rect 35156 37562 35180 37564
rect 35236 37562 35242 37564
rect 34996 37510 34998 37562
rect 35178 37510 35180 37562
rect 34934 37508 34940 37510
rect 34996 37508 35020 37510
rect 35076 37508 35100 37510
rect 35156 37508 35180 37510
rect 35236 37508 35242 37510
rect 34934 37488 35242 37508
rect 34934 36476 35242 36496
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36400 35242 36420
rect 34934 35388 35242 35408
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35312 35242 35332
rect 34934 34300 35242 34320
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34224 35242 34244
rect 34934 33212 35242 33232
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33136 35242 33156
rect 34934 32124 35242 32144
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32048 35242 32068
rect 34934 31036 35242 31056
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30960 35242 30980
rect 34934 29948 35242 29968
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29872 35242 29892
rect 34934 28860 35242 28880
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28784 35242 28804
rect 34934 27772 35242 27792
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27696 35242 27716
rect 34934 26684 35242 26704
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26608 35242 26628
rect 34934 25596 35242 25616
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25520 35242 25540
rect 34934 24508 35242 24528
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24432 35242 24452
rect 34934 23420 35242 23440
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23344 35242 23364
rect 34934 22332 35242 22352
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22256 35242 22276
rect 34934 21244 35242 21264
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21168 35242 21188
rect 34934 20156 35242 20176
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20080 35242 20100
rect 34934 19068 35242 19088
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 18992 35242 19012
rect 34934 17980 35242 18000
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17904 35242 17924
rect 34934 16892 35242 16912
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16816 35242 16836
rect 34934 15804 35242 15824
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15728 35242 15748
rect 34934 14716 35242 14736
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14640 35242 14660
rect 34934 13628 35242 13648
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13552 35242 13572
rect 34934 12540 35242 12560
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12464 35242 12484
rect 34934 11452 35242 11472
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11376 35242 11396
rect 34934 10364 35242 10384
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10288 35242 10308
rect 34934 9276 35242 9296
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9200 35242 9220
rect 34934 8188 35242 8208
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8112 35242 8132
rect 34934 7100 35242 7120
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7024 35242 7044
rect 34934 6012 35242 6032
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5936 35242 5956
rect 34934 4924 35242 4944
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4848 35242 4868
rect 34934 3836 35242 3856
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3760 35242 3780
rect 34934 2748 35242 2768
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2672 35242 2692
rect 29920 2644 29972 2650
rect 29920 2586 29972 2592
rect 33140 2644 33192 2650
rect 33140 2586 33192 2592
rect 19984 2508 20036 2514
rect 19984 2450 20036 2456
rect 35360 2446 35388 59910
rect 36280 59770 36308 59978
rect 37740 59968 37792 59974
rect 37740 59910 37792 59916
rect 36268 59764 36320 59770
rect 36268 59706 36320 59712
rect 37752 59702 37780 59910
rect 37740 59696 37792 59702
rect 37740 59638 37792 59644
rect 38856 38758 38884 60658
rect 38936 60036 38988 60042
rect 38936 59978 38988 59984
rect 38844 38752 38896 38758
rect 38844 38694 38896 38700
rect 38948 23662 38976 59978
rect 39120 59560 39172 59566
rect 39120 59502 39172 59508
rect 39132 24614 39160 59502
rect 39500 50930 39528 63718
rect 39764 61192 39816 61198
rect 39764 61134 39816 61140
rect 39580 59628 39632 59634
rect 39580 59570 39632 59576
rect 39488 50924 39540 50930
rect 39488 50866 39540 50872
rect 39592 43110 39620 59570
rect 39672 59016 39724 59022
rect 39672 58958 39724 58964
rect 39580 43104 39632 43110
rect 39580 43046 39632 43052
rect 39684 27402 39712 58958
rect 39672 27396 39724 27402
rect 39672 27338 39724 27344
rect 39580 25696 39632 25702
rect 39580 25638 39632 25644
rect 39592 25498 39620 25638
rect 39580 25492 39632 25498
rect 39580 25434 39632 25440
rect 39120 24608 39172 24614
rect 39120 24550 39172 24556
rect 38936 23656 38988 23662
rect 38936 23598 38988 23604
rect 3240 2440 3292 2446
rect 3240 2382 3292 2388
rect 7104 2440 7156 2446
rect 7104 2382 7156 2388
rect 11520 2440 11572 2446
rect 11520 2382 11572 2388
rect 16212 2440 16264 2446
rect 16212 2382 16264 2388
rect 29644 2440 29696 2446
rect 29644 2382 29696 2388
rect 35348 2440 35400 2446
rect 35348 2382 35400 2388
rect 2964 2032 3016 2038
rect 2964 1974 3016 1980
rect 3252 800 3280 2382
rect 7116 800 7144 2382
rect 7840 2372 7892 2378
rect 7840 2314 7892 2320
rect 14832 2372 14884 2378
rect 14832 2314 14884 2320
rect 18052 2372 18104 2378
rect 18052 2314 18104 2320
rect 7852 1902 7880 2314
rect 10968 2304 11020 2310
rect 10968 2246 11020 2252
rect 7840 1896 7892 1902
rect 7840 1838 7892 1844
rect 10980 800 11008 2246
rect 14844 800 14872 2314
rect 18064 800 18092 2314
rect 21916 2304 21968 2310
rect 21916 2246 21968 2252
rect 25780 2304 25832 2310
rect 25780 2246 25832 2252
rect 19574 2204 19882 2224
rect 19574 2202 19580 2204
rect 19636 2202 19660 2204
rect 19716 2202 19740 2204
rect 19796 2202 19820 2204
rect 19876 2202 19882 2204
rect 19636 2150 19638 2202
rect 19818 2150 19820 2202
rect 19574 2148 19580 2150
rect 19636 2148 19660 2150
rect 19716 2148 19740 2150
rect 19796 2148 19820 2150
rect 19876 2148 19882 2150
rect 19574 2128 19882 2148
rect 21928 800 21956 2246
rect 25792 800 25820 2246
rect 29656 800 29684 2382
rect 39776 2378 39804 61134
rect 39868 48278 39896 65486
rect 40040 65476 40092 65482
rect 40040 65418 40092 65424
rect 40052 65210 40080 65418
rect 40040 65204 40092 65210
rect 40040 65146 40092 65152
rect 40696 65006 40724 65554
rect 41064 65210 41092 89966
rect 45204 72010 45232 117234
rect 45388 117162 45416 119326
rect 48962 119326 49280 119354
rect 48962 119200 49018 119326
rect 49252 117298 49280 119326
rect 52182 119326 52408 119354
rect 52182 119200 52238 119326
rect 50294 117532 50602 117552
rect 50294 117530 50300 117532
rect 50356 117530 50380 117532
rect 50436 117530 50460 117532
rect 50516 117530 50540 117532
rect 50596 117530 50602 117532
rect 50356 117478 50358 117530
rect 50538 117478 50540 117530
rect 50294 117476 50300 117478
rect 50356 117476 50380 117478
rect 50436 117476 50460 117478
rect 50516 117476 50540 117478
rect 50596 117476 50602 117478
rect 50294 117456 50602 117476
rect 49240 117292 49292 117298
rect 49240 117234 49292 117240
rect 45376 117156 45428 117162
rect 52380 117144 52408 119326
rect 56046 119326 56180 119354
rect 56046 119200 56102 119326
rect 56152 117298 56180 119326
rect 59910 119200 59966 120000
rect 63774 119354 63830 120000
rect 66994 119354 67050 120000
rect 63774 119326 64092 119354
rect 63774 119200 63830 119326
rect 59924 117298 59952 119200
rect 56140 117292 56192 117298
rect 56140 117234 56192 117240
rect 59912 117292 59964 117298
rect 59912 117234 59964 117240
rect 63868 117292 63920 117298
rect 63868 117234 63920 117240
rect 56324 117224 56376 117230
rect 56324 117166 56376 117172
rect 52460 117156 52512 117162
rect 52380 117116 52460 117144
rect 45376 117098 45428 117104
rect 52460 117098 52512 117104
rect 49056 117088 49108 117094
rect 49056 117030 49108 117036
rect 49068 116210 49096 117030
rect 50294 116444 50602 116464
rect 50294 116442 50300 116444
rect 50356 116442 50380 116444
rect 50436 116442 50460 116444
rect 50516 116442 50540 116444
rect 50596 116442 50602 116444
rect 50356 116390 50358 116442
rect 50538 116390 50540 116442
rect 50294 116388 50300 116390
rect 50356 116388 50380 116390
rect 50436 116388 50460 116390
rect 50516 116388 50540 116390
rect 50596 116388 50602 116390
rect 50294 116368 50602 116388
rect 49056 116204 49108 116210
rect 49056 116146 49108 116152
rect 50294 115356 50602 115376
rect 50294 115354 50300 115356
rect 50356 115354 50380 115356
rect 50436 115354 50460 115356
rect 50516 115354 50540 115356
rect 50596 115354 50602 115356
rect 50356 115302 50358 115354
rect 50538 115302 50540 115354
rect 50294 115300 50300 115302
rect 50356 115300 50380 115302
rect 50436 115300 50460 115302
rect 50516 115300 50540 115302
rect 50596 115300 50602 115302
rect 50294 115280 50602 115300
rect 50294 114268 50602 114288
rect 50294 114266 50300 114268
rect 50356 114266 50380 114268
rect 50436 114266 50460 114268
rect 50516 114266 50540 114268
rect 50596 114266 50602 114268
rect 50356 114214 50358 114266
rect 50538 114214 50540 114266
rect 50294 114212 50300 114214
rect 50356 114212 50380 114214
rect 50436 114212 50460 114214
rect 50516 114212 50540 114214
rect 50596 114212 50602 114214
rect 50294 114192 50602 114212
rect 50294 113180 50602 113200
rect 50294 113178 50300 113180
rect 50356 113178 50380 113180
rect 50436 113178 50460 113180
rect 50516 113178 50540 113180
rect 50596 113178 50602 113180
rect 50356 113126 50358 113178
rect 50538 113126 50540 113178
rect 50294 113124 50300 113126
rect 50356 113124 50380 113126
rect 50436 113124 50460 113126
rect 50516 113124 50540 113126
rect 50596 113124 50602 113126
rect 50294 113104 50602 113124
rect 50294 112092 50602 112112
rect 50294 112090 50300 112092
rect 50356 112090 50380 112092
rect 50436 112090 50460 112092
rect 50516 112090 50540 112092
rect 50596 112090 50602 112092
rect 50356 112038 50358 112090
rect 50538 112038 50540 112090
rect 50294 112036 50300 112038
rect 50356 112036 50380 112038
rect 50436 112036 50460 112038
rect 50516 112036 50540 112038
rect 50596 112036 50602 112038
rect 50294 112016 50602 112036
rect 50294 111004 50602 111024
rect 50294 111002 50300 111004
rect 50356 111002 50380 111004
rect 50436 111002 50460 111004
rect 50516 111002 50540 111004
rect 50596 111002 50602 111004
rect 50356 110950 50358 111002
rect 50538 110950 50540 111002
rect 50294 110948 50300 110950
rect 50356 110948 50380 110950
rect 50436 110948 50460 110950
rect 50516 110948 50540 110950
rect 50596 110948 50602 110950
rect 50294 110928 50602 110948
rect 50294 109916 50602 109936
rect 50294 109914 50300 109916
rect 50356 109914 50380 109916
rect 50436 109914 50460 109916
rect 50516 109914 50540 109916
rect 50596 109914 50602 109916
rect 50356 109862 50358 109914
rect 50538 109862 50540 109914
rect 50294 109860 50300 109862
rect 50356 109860 50380 109862
rect 50436 109860 50460 109862
rect 50516 109860 50540 109862
rect 50596 109860 50602 109862
rect 50294 109840 50602 109860
rect 50294 108828 50602 108848
rect 50294 108826 50300 108828
rect 50356 108826 50380 108828
rect 50436 108826 50460 108828
rect 50516 108826 50540 108828
rect 50596 108826 50602 108828
rect 50356 108774 50358 108826
rect 50538 108774 50540 108826
rect 50294 108772 50300 108774
rect 50356 108772 50380 108774
rect 50436 108772 50460 108774
rect 50516 108772 50540 108774
rect 50596 108772 50602 108774
rect 50294 108752 50602 108772
rect 50294 107740 50602 107760
rect 50294 107738 50300 107740
rect 50356 107738 50380 107740
rect 50436 107738 50460 107740
rect 50516 107738 50540 107740
rect 50596 107738 50602 107740
rect 50356 107686 50358 107738
rect 50538 107686 50540 107738
rect 50294 107684 50300 107686
rect 50356 107684 50380 107686
rect 50436 107684 50460 107686
rect 50516 107684 50540 107686
rect 50596 107684 50602 107686
rect 50294 107664 50602 107684
rect 50294 106652 50602 106672
rect 50294 106650 50300 106652
rect 50356 106650 50380 106652
rect 50436 106650 50460 106652
rect 50516 106650 50540 106652
rect 50596 106650 50602 106652
rect 50356 106598 50358 106650
rect 50538 106598 50540 106650
rect 50294 106596 50300 106598
rect 50356 106596 50380 106598
rect 50436 106596 50460 106598
rect 50516 106596 50540 106598
rect 50596 106596 50602 106598
rect 50294 106576 50602 106596
rect 50294 105564 50602 105584
rect 50294 105562 50300 105564
rect 50356 105562 50380 105564
rect 50436 105562 50460 105564
rect 50516 105562 50540 105564
rect 50596 105562 50602 105564
rect 50356 105510 50358 105562
rect 50538 105510 50540 105562
rect 50294 105508 50300 105510
rect 50356 105508 50380 105510
rect 50436 105508 50460 105510
rect 50516 105508 50540 105510
rect 50596 105508 50602 105510
rect 50294 105488 50602 105508
rect 50294 104476 50602 104496
rect 50294 104474 50300 104476
rect 50356 104474 50380 104476
rect 50436 104474 50460 104476
rect 50516 104474 50540 104476
rect 50596 104474 50602 104476
rect 50356 104422 50358 104474
rect 50538 104422 50540 104474
rect 50294 104420 50300 104422
rect 50356 104420 50380 104422
rect 50436 104420 50460 104422
rect 50516 104420 50540 104422
rect 50596 104420 50602 104422
rect 50294 104400 50602 104420
rect 50294 103388 50602 103408
rect 50294 103386 50300 103388
rect 50356 103386 50380 103388
rect 50436 103386 50460 103388
rect 50516 103386 50540 103388
rect 50596 103386 50602 103388
rect 50356 103334 50358 103386
rect 50538 103334 50540 103386
rect 50294 103332 50300 103334
rect 50356 103332 50380 103334
rect 50436 103332 50460 103334
rect 50516 103332 50540 103334
rect 50596 103332 50602 103334
rect 50294 103312 50602 103332
rect 50294 102300 50602 102320
rect 50294 102298 50300 102300
rect 50356 102298 50380 102300
rect 50436 102298 50460 102300
rect 50516 102298 50540 102300
rect 50596 102298 50602 102300
rect 50356 102246 50358 102298
rect 50538 102246 50540 102298
rect 50294 102244 50300 102246
rect 50356 102244 50380 102246
rect 50436 102244 50460 102246
rect 50516 102244 50540 102246
rect 50596 102244 50602 102246
rect 50294 102224 50602 102244
rect 50294 101212 50602 101232
rect 50294 101210 50300 101212
rect 50356 101210 50380 101212
rect 50436 101210 50460 101212
rect 50516 101210 50540 101212
rect 50596 101210 50602 101212
rect 50356 101158 50358 101210
rect 50538 101158 50540 101210
rect 50294 101156 50300 101158
rect 50356 101156 50380 101158
rect 50436 101156 50460 101158
rect 50516 101156 50540 101158
rect 50596 101156 50602 101158
rect 50294 101136 50602 101156
rect 50294 100124 50602 100144
rect 50294 100122 50300 100124
rect 50356 100122 50380 100124
rect 50436 100122 50460 100124
rect 50516 100122 50540 100124
rect 50596 100122 50602 100124
rect 50356 100070 50358 100122
rect 50538 100070 50540 100122
rect 50294 100068 50300 100070
rect 50356 100068 50380 100070
rect 50436 100068 50460 100070
rect 50516 100068 50540 100070
rect 50596 100068 50602 100070
rect 50294 100048 50602 100068
rect 50294 99036 50602 99056
rect 50294 99034 50300 99036
rect 50356 99034 50380 99036
rect 50436 99034 50460 99036
rect 50516 99034 50540 99036
rect 50596 99034 50602 99036
rect 50356 98982 50358 99034
rect 50538 98982 50540 99034
rect 50294 98980 50300 98982
rect 50356 98980 50380 98982
rect 50436 98980 50460 98982
rect 50516 98980 50540 98982
rect 50596 98980 50602 98982
rect 50294 98960 50602 98980
rect 50294 97948 50602 97968
rect 50294 97946 50300 97948
rect 50356 97946 50380 97948
rect 50436 97946 50460 97948
rect 50516 97946 50540 97948
rect 50596 97946 50602 97948
rect 50356 97894 50358 97946
rect 50538 97894 50540 97946
rect 50294 97892 50300 97894
rect 50356 97892 50380 97894
rect 50436 97892 50460 97894
rect 50516 97892 50540 97894
rect 50596 97892 50602 97894
rect 50294 97872 50602 97892
rect 50294 96860 50602 96880
rect 50294 96858 50300 96860
rect 50356 96858 50380 96860
rect 50436 96858 50460 96860
rect 50516 96858 50540 96860
rect 50596 96858 50602 96860
rect 50356 96806 50358 96858
rect 50538 96806 50540 96858
rect 50294 96804 50300 96806
rect 50356 96804 50380 96806
rect 50436 96804 50460 96806
rect 50516 96804 50540 96806
rect 50596 96804 50602 96806
rect 50294 96784 50602 96804
rect 50294 95772 50602 95792
rect 50294 95770 50300 95772
rect 50356 95770 50380 95772
rect 50436 95770 50460 95772
rect 50516 95770 50540 95772
rect 50596 95770 50602 95772
rect 50356 95718 50358 95770
rect 50538 95718 50540 95770
rect 50294 95716 50300 95718
rect 50356 95716 50380 95718
rect 50436 95716 50460 95718
rect 50516 95716 50540 95718
rect 50596 95716 50602 95718
rect 50294 95696 50602 95716
rect 50294 94684 50602 94704
rect 50294 94682 50300 94684
rect 50356 94682 50380 94684
rect 50436 94682 50460 94684
rect 50516 94682 50540 94684
rect 50596 94682 50602 94684
rect 50356 94630 50358 94682
rect 50538 94630 50540 94682
rect 50294 94628 50300 94630
rect 50356 94628 50380 94630
rect 50436 94628 50460 94630
rect 50516 94628 50540 94630
rect 50596 94628 50602 94630
rect 50294 94608 50602 94628
rect 50294 93596 50602 93616
rect 50294 93594 50300 93596
rect 50356 93594 50380 93596
rect 50436 93594 50460 93596
rect 50516 93594 50540 93596
rect 50596 93594 50602 93596
rect 50356 93542 50358 93594
rect 50538 93542 50540 93594
rect 50294 93540 50300 93542
rect 50356 93540 50380 93542
rect 50436 93540 50460 93542
rect 50516 93540 50540 93542
rect 50596 93540 50602 93542
rect 50294 93520 50602 93540
rect 50294 92508 50602 92528
rect 50294 92506 50300 92508
rect 50356 92506 50380 92508
rect 50436 92506 50460 92508
rect 50516 92506 50540 92508
rect 50596 92506 50602 92508
rect 50356 92454 50358 92506
rect 50538 92454 50540 92506
rect 50294 92452 50300 92454
rect 50356 92452 50380 92454
rect 50436 92452 50460 92454
rect 50516 92452 50540 92454
rect 50596 92452 50602 92454
rect 50294 92432 50602 92452
rect 50294 91420 50602 91440
rect 50294 91418 50300 91420
rect 50356 91418 50380 91420
rect 50436 91418 50460 91420
rect 50516 91418 50540 91420
rect 50596 91418 50602 91420
rect 50356 91366 50358 91418
rect 50538 91366 50540 91418
rect 50294 91364 50300 91366
rect 50356 91364 50380 91366
rect 50436 91364 50460 91366
rect 50516 91364 50540 91366
rect 50596 91364 50602 91366
rect 50294 91344 50602 91364
rect 50294 90332 50602 90352
rect 50294 90330 50300 90332
rect 50356 90330 50380 90332
rect 50436 90330 50460 90332
rect 50516 90330 50540 90332
rect 50596 90330 50602 90332
rect 50356 90278 50358 90330
rect 50538 90278 50540 90330
rect 50294 90276 50300 90278
rect 50356 90276 50380 90278
rect 50436 90276 50460 90278
rect 50516 90276 50540 90278
rect 50596 90276 50602 90278
rect 50294 90256 50602 90276
rect 50294 89244 50602 89264
rect 50294 89242 50300 89244
rect 50356 89242 50380 89244
rect 50436 89242 50460 89244
rect 50516 89242 50540 89244
rect 50596 89242 50602 89244
rect 50356 89190 50358 89242
rect 50538 89190 50540 89242
rect 50294 89188 50300 89190
rect 50356 89188 50380 89190
rect 50436 89188 50460 89190
rect 50516 89188 50540 89190
rect 50596 89188 50602 89190
rect 50294 89168 50602 89188
rect 50294 88156 50602 88176
rect 50294 88154 50300 88156
rect 50356 88154 50380 88156
rect 50436 88154 50460 88156
rect 50516 88154 50540 88156
rect 50596 88154 50602 88156
rect 50356 88102 50358 88154
rect 50538 88102 50540 88154
rect 50294 88100 50300 88102
rect 50356 88100 50380 88102
rect 50436 88100 50460 88102
rect 50516 88100 50540 88102
rect 50596 88100 50602 88102
rect 50294 88080 50602 88100
rect 50294 87068 50602 87088
rect 50294 87066 50300 87068
rect 50356 87066 50380 87068
rect 50436 87066 50460 87068
rect 50516 87066 50540 87068
rect 50596 87066 50602 87068
rect 50356 87014 50358 87066
rect 50538 87014 50540 87066
rect 50294 87012 50300 87014
rect 50356 87012 50380 87014
rect 50436 87012 50460 87014
rect 50516 87012 50540 87014
rect 50596 87012 50602 87014
rect 50294 86992 50602 87012
rect 50294 85980 50602 86000
rect 50294 85978 50300 85980
rect 50356 85978 50380 85980
rect 50436 85978 50460 85980
rect 50516 85978 50540 85980
rect 50596 85978 50602 85980
rect 50356 85926 50358 85978
rect 50538 85926 50540 85978
rect 50294 85924 50300 85926
rect 50356 85924 50380 85926
rect 50436 85924 50460 85926
rect 50516 85924 50540 85926
rect 50596 85924 50602 85926
rect 50294 85904 50602 85924
rect 50294 84892 50602 84912
rect 50294 84890 50300 84892
rect 50356 84890 50380 84892
rect 50436 84890 50460 84892
rect 50516 84890 50540 84892
rect 50596 84890 50602 84892
rect 50356 84838 50358 84890
rect 50538 84838 50540 84890
rect 50294 84836 50300 84838
rect 50356 84836 50380 84838
rect 50436 84836 50460 84838
rect 50516 84836 50540 84838
rect 50596 84836 50602 84838
rect 50294 84816 50602 84836
rect 50294 83804 50602 83824
rect 50294 83802 50300 83804
rect 50356 83802 50380 83804
rect 50436 83802 50460 83804
rect 50516 83802 50540 83804
rect 50596 83802 50602 83804
rect 50356 83750 50358 83802
rect 50538 83750 50540 83802
rect 50294 83748 50300 83750
rect 50356 83748 50380 83750
rect 50436 83748 50460 83750
rect 50516 83748 50540 83750
rect 50596 83748 50602 83750
rect 50294 83728 50602 83748
rect 50294 82716 50602 82736
rect 50294 82714 50300 82716
rect 50356 82714 50380 82716
rect 50436 82714 50460 82716
rect 50516 82714 50540 82716
rect 50596 82714 50602 82716
rect 50356 82662 50358 82714
rect 50538 82662 50540 82714
rect 50294 82660 50300 82662
rect 50356 82660 50380 82662
rect 50436 82660 50460 82662
rect 50516 82660 50540 82662
rect 50596 82660 50602 82662
rect 50294 82640 50602 82660
rect 50294 81628 50602 81648
rect 50294 81626 50300 81628
rect 50356 81626 50380 81628
rect 50436 81626 50460 81628
rect 50516 81626 50540 81628
rect 50596 81626 50602 81628
rect 50356 81574 50358 81626
rect 50538 81574 50540 81626
rect 50294 81572 50300 81574
rect 50356 81572 50380 81574
rect 50436 81572 50460 81574
rect 50516 81572 50540 81574
rect 50596 81572 50602 81574
rect 50294 81552 50602 81572
rect 50294 80540 50602 80560
rect 50294 80538 50300 80540
rect 50356 80538 50380 80540
rect 50436 80538 50460 80540
rect 50516 80538 50540 80540
rect 50596 80538 50602 80540
rect 50356 80486 50358 80538
rect 50538 80486 50540 80538
rect 50294 80484 50300 80486
rect 50356 80484 50380 80486
rect 50436 80484 50460 80486
rect 50516 80484 50540 80486
rect 50596 80484 50602 80486
rect 50294 80464 50602 80484
rect 50294 79452 50602 79472
rect 50294 79450 50300 79452
rect 50356 79450 50380 79452
rect 50436 79450 50460 79452
rect 50516 79450 50540 79452
rect 50596 79450 50602 79452
rect 50356 79398 50358 79450
rect 50538 79398 50540 79450
rect 50294 79396 50300 79398
rect 50356 79396 50380 79398
rect 50436 79396 50460 79398
rect 50516 79396 50540 79398
rect 50596 79396 50602 79398
rect 50294 79376 50602 79396
rect 50294 78364 50602 78384
rect 50294 78362 50300 78364
rect 50356 78362 50380 78364
rect 50436 78362 50460 78364
rect 50516 78362 50540 78364
rect 50596 78362 50602 78364
rect 50356 78310 50358 78362
rect 50538 78310 50540 78362
rect 50294 78308 50300 78310
rect 50356 78308 50380 78310
rect 50436 78308 50460 78310
rect 50516 78308 50540 78310
rect 50596 78308 50602 78310
rect 50294 78288 50602 78308
rect 50294 77276 50602 77296
rect 50294 77274 50300 77276
rect 50356 77274 50380 77276
rect 50436 77274 50460 77276
rect 50516 77274 50540 77276
rect 50596 77274 50602 77276
rect 50356 77222 50358 77274
rect 50538 77222 50540 77274
rect 50294 77220 50300 77222
rect 50356 77220 50380 77222
rect 50436 77220 50460 77222
rect 50516 77220 50540 77222
rect 50596 77220 50602 77222
rect 50294 77200 50602 77220
rect 50294 76188 50602 76208
rect 50294 76186 50300 76188
rect 50356 76186 50380 76188
rect 50436 76186 50460 76188
rect 50516 76186 50540 76188
rect 50596 76186 50602 76188
rect 50356 76134 50358 76186
rect 50538 76134 50540 76186
rect 50294 76132 50300 76134
rect 50356 76132 50380 76134
rect 50436 76132 50460 76134
rect 50516 76132 50540 76134
rect 50596 76132 50602 76134
rect 50294 76112 50602 76132
rect 50294 75100 50602 75120
rect 50294 75098 50300 75100
rect 50356 75098 50380 75100
rect 50436 75098 50460 75100
rect 50516 75098 50540 75100
rect 50596 75098 50602 75100
rect 50356 75046 50358 75098
rect 50538 75046 50540 75098
rect 50294 75044 50300 75046
rect 50356 75044 50380 75046
rect 50436 75044 50460 75046
rect 50516 75044 50540 75046
rect 50596 75044 50602 75046
rect 50294 75024 50602 75044
rect 50294 74012 50602 74032
rect 50294 74010 50300 74012
rect 50356 74010 50380 74012
rect 50436 74010 50460 74012
rect 50516 74010 50540 74012
rect 50596 74010 50602 74012
rect 50356 73958 50358 74010
rect 50538 73958 50540 74010
rect 50294 73956 50300 73958
rect 50356 73956 50380 73958
rect 50436 73956 50460 73958
rect 50516 73956 50540 73958
rect 50596 73956 50602 73958
rect 50294 73936 50602 73956
rect 50294 72924 50602 72944
rect 50294 72922 50300 72924
rect 50356 72922 50380 72924
rect 50436 72922 50460 72924
rect 50516 72922 50540 72924
rect 50596 72922 50602 72924
rect 50356 72870 50358 72922
rect 50538 72870 50540 72922
rect 50294 72868 50300 72870
rect 50356 72868 50380 72870
rect 50436 72868 50460 72870
rect 50516 72868 50540 72870
rect 50596 72868 50602 72870
rect 50294 72848 50602 72868
rect 45192 72004 45244 72010
rect 45192 71946 45244 71952
rect 50294 71836 50602 71856
rect 50294 71834 50300 71836
rect 50356 71834 50380 71836
rect 50436 71834 50460 71836
rect 50516 71834 50540 71836
rect 50596 71834 50602 71836
rect 50356 71782 50358 71834
rect 50538 71782 50540 71834
rect 50294 71780 50300 71782
rect 50356 71780 50380 71782
rect 50436 71780 50460 71782
rect 50516 71780 50540 71782
rect 50596 71780 50602 71782
rect 50294 71760 50602 71780
rect 50294 70748 50602 70768
rect 50294 70746 50300 70748
rect 50356 70746 50380 70748
rect 50436 70746 50460 70748
rect 50516 70746 50540 70748
rect 50596 70746 50602 70748
rect 50356 70694 50358 70746
rect 50538 70694 50540 70746
rect 50294 70692 50300 70694
rect 50356 70692 50380 70694
rect 50436 70692 50460 70694
rect 50516 70692 50540 70694
rect 50596 70692 50602 70694
rect 50294 70672 50602 70692
rect 50294 69660 50602 69680
rect 50294 69658 50300 69660
rect 50356 69658 50380 69660
rect 50436 69658 50460 69660
rect 50516 69658 50540 69660
rect 50596 69658 50602 69660
rect 50356 69606 50358 69658
rect 50538 69606 50540 69658
rect 50294 69604 50300 69606
rect 50356 69604 50380 69606
rect 50436 69604 50460 69606
rect 50516 69604 50540 69606
rect 50596 69604 50602 69606
rect 50294 69584 50602 69604
rect 50294 68572 50602 68592
rect 50294 68570 50300 68572
rect 50356 68570 50380 68572
rect 50436 68570 50460 68572
rect 50516 68570 50540 68572
rect 50596 68570 50602 68572
rect 50356 68518 50358 68570
rect 50538 68518 50540 68570
rect 50294 68516 50300 68518
rect 50356 68516 50380 68518
rect 50436 68516 50460 68518
rect 50516 68516 50540 68518
rect 50596 68516 50602 68518
rect 50294 68496 50602 68516
rect 50294 67484 50602 67504
rect 50294 67482 50300 67484
rect 50356 67482 50380 67484
rect 50436 67482 50460 67484
rect 50516 67482 50540 67484
rect 50596 67482 50602 67484
rect 50356 67430 50358 67482
rect 50538 67430 50540 67482
rect 50294 67428 50300 67430
rect 50356 67428 50380 67430
rect 50436 67428 50460 67430
rect 50516 67428 50540 67430
rect 50596 67428 50602 67430
rect 50294 67408 50602 67428
rect 50294 66396 50602 66416
rect 50294 66394 50300 66396
rect 50356 66394 50380 66396
rect 50436 66394 50460 66396
rect 50516 66394 50540 66396
rect 50596 66394 50602 66396
rect 50356 66342 50358 66394
rect 50538 66342 50540 66394
rect 50294 66340 50300 66342
rect 50356 66340 50380 66342
rect 50436 66340 50460 66342
rect 50516 66340 50540 66342
rect 50596 66340 50602 66342
rect 50294 66320 50602 66340
rect 50294 65308 50602 65328
rect 50294 65306 50300 65308
rect 50356 65306 50380 65308
rect 50436 65306 50460 65308
rect 50516 65306 50540 65308
rect 50596 65306 50602 65308
rect 50356 65254 50358 65306
rect 50538 65254 50540 65306
rect 50294 65252 50300 65254
rect 50356 65252 50380 65254
rect 50436 65252 50460 65254
rect 50516 65252 50540 65254
rect 50596 65252 50602 65254
rect 50294 65232 50602 65252
rect 41052 65204 41104 65210
rect 41052 65146 41104 65152
rect 40684 65000 40736 65006
rect 40684 64942 40736 64948
rect 40868 64864 40920 64870
rect 40868 64806 40920 64812
rect 40880 64462 40908 64806
rect 41064 64530 41092 65146
rect 41696 64864 41748 64870
rect 41696 64806 41748 64812
rect 41708 64598 41736 64806
rect 41696 64592 41748 64598
rect 41696 64534 41748 64540
rect 41052 64524 41104 64530
rect 41052 64466 41104 64472
rect 40500 64456 40552 64462
rect 40500 64398 40552 64404
rect 40868 64456 40920 64462
rect 40868 64398 40920 64404
rect 39948 60784 40000 60790
rect 39948 60726 40000 60732
rect 39856 48272 39908 48278
rect 39856 48214 39908 48220
rect 32864 2372 32916 2378
rect 32864 2314 32916 2320
rect 39764 2372 39816 2378
rect 39764 2314 39816 2320
rect 32876 800 32904 2314
rect 36728 2304 36780 2310
rect 36728 2246 36780 2252
rect 36740 800 36768 2246
rect 39960 1970 39988 60726
rect 40512 54670 40540 64398
rect 40776 60784 40828 60790
rect 40776 60726 40828 60732
rect 40592 60036 40644 60042
rect 40592 59978 40644 59984
rect 40500 54664 40552 54670
rect 40500 54606 40552 54612
rect 40604 8838 40632 59978
rect 40788 31890 40816 60726
rect 40776 31884 40828 31890
rect 40776 31826 40828 31832
rect 40592 8832 40644 8838
rect 40592 8774 40644 8780
rect 40408 3392 40460 3398
rect 40408 3334 40460 3340
rect 40420 3194 40448 3334
rect 40408 3188 40460 3194
rect 40408 3130 40460 3136
rect 40880 2530 40908 64398
rect 50294 64220 50602 64240
rect 50294 64218 50300 64220
rect 50356 64218 50380 64220
rect 50436 64218 50460 64220
rect 50516 64218 50540 64220
rect 50596 64218 50602 64220
rect 50356 64166 50358 64218
rect 50538 64166 50540 64218
rect 50294 64164 50300 64166
rect 50356 64164 50380 64166
rect 50436 64164 50460 64166
rect 50516 64164 50540 64166
rect 50596 64164 50602 64166
rect 50294 64144 50602 64164
rect 50294 63132 50602 63152
rect 50294 63130 50300 63132
rect 50356 63130 50380 63132
rect 50436 63130 50460 63132
rect 50516 63130 50540 63132
rect 50596 63130 50602 63132
rect 50356 63078 50358 63130
rect 50538 63078 50540 63130
rect 50294 63076 50300 63078
rect 50356 63076 50380 63078
rect 50436 63076 50460 63078
rect 50516 63076 50540 63078
rect 50596 63076 50602 63078
rect 50294 63056 50602 63076
rect 50294 62044 50602 62064
rect 50294 62042 50300 62044
rect 50356 62042 50380 62044
rect 50436 62042 50460 62044
rect 50516 62042 50540 62044
rect 50596 62042 50602 62044
rect 50356 61990 50358 62042
rect 50538 61990 50540 62042
rect 50294 61988 50300 61990
rect 50356 61988 50380 61990
rect 50436 61988 50460 61990
rect 50516 61988 50540 61990
rect 50596 61988 50602 61990
rect 50294 61968 50602 61988
rect 50294 60956 50602 60976
rect 50294 60954 50300 60956
rect 50356 60954 50380 60956
rect 50436 60954 50460 60956
rect 50516 60954 50540 60956
rect 50596 60954 50602 60956
rect 50356 60902 50358 60954
rect 50538 60902 50540 60954
rect 50294 60900 50300 60902
rect 50356 60900 50380 60902
rect 50436 60900 50460 60902
rect 50516 60900 50540 60902
rect 50596 60900 50602 60902
rect 50294 60880 50602 60900
rect 56336 60110 56364 117166
rect 58624 117156 58676 117162
rect 58624 117098 58676 117104
rect 58636 100570 58664 117098
rect 58624 100564 58676 100570
rect 58624 100506 58676 100512
rect 58532 100292 58584 100298
rect 58532 100234 58584 100240
rect 58544 90438 58572 100234
rect 58532 90432 58584 90438
rect 58532 90374 58584 90380
rect 41052 60104 41104 60110
rect 41052 60046 41104 60052
rect 56324 60104 56376 60110
rect 56324 60046 56376 60052
rect 40960 3528 41012 3534
rect 40960 3470 41012 3476
rect 40972 2650 41000 3470
rect 40960 2644 41012 2650
rect 40960 2586 41012 2592
rect 41064 2582 41092 60046
rect 63040 59968 63092 59974
rect 63040 59910 63092 59916
rect 50294 59868 50602 59888
rect 50294 59866 50300 59868
rect 50356 59866 50380 59868
rect 50436 59866 50460 59868
rect 50516 59866 50540 59868
rect 50596 59866 50602 59868
rect 50356 59814 50358 59866
rect 50538 59814 50540 59866
rect 50294 59812 50300 59814
rect 50356 59812 50380 59814
rect 50436 59812 50460 59814
rect 50516 59812 50540 59814
rect 50596 59812 50602 59814
rect 50294 59792 50602 59812
rect 41144 59628 41196 59634
rect 41144 59570 41196 59576
rect 41156 16574 41184 59570
rect 50294 58780 50602 58800
rect 50294 58778 50300 58780
rect 50356 58778 50380 58780
rect 50436 58778 50460 58780
rect 50516 58778 50540 58780
rect 50596 58778 50602 58780
rect 50356 58726 50358 58778
rect 50538 58726 50540 58778
rect 50294 58724 50300 58726
rect 50356 58724 50380 58726
rect 50436 58724 50460 58726
rect 50516 58724 50540 58726
rect 50596 58724 50602 58726
rect 50294 58704 50602 58724
rect 50294 57692 50602 57712
rect 50294 57690 50300 57692
rect 50356 57690 50380 57692
rect 50436 57690 50460 57692
rect 50516 57690 50540 57692
rect 50596 57690 50602 57692
rect 50356 57638 50358 57690
rect 50538 57638 50540 57690
rect 50294 57636 50300 57638
rect 50356 57636 50380 57638
rect 50436 57636 50460 57638
rect 50516 57636 50540 57638
rect 50596 57636 50602 57638
rect 50294 57616 50602 57636
rect 50294 56604 50602 56624
rect 50294 56602 50300 56604
rect 50356 56602 50380 56604
rect 50436 56602 50460 56604
rect 50516 56602 50540 56604
rect 50596 56602 50602 56604
rect 50356 56550 50358 56602
rect 50538 56550 50540 56602
rect 50294 56548 50300 56550
rect 50356 56548 50380 56550
rect 50436 56548 50460 56550
rect 50516 56548 50540 56550
rect 50596 56548 50602 56550
rect 50294 56528 50602 56548
rect 50294 55516 50602 55536
rect 50294 55514 50300 55516
rect 50356 55514 50380 55516
rect 50436 55514 50460 55516
rect 50516 55514 50540 55516
rect 50596 55514 50602 55516
rect 50356 55462 50358 55514
rect 50538 55462 50540 55514
rect 50294 55460 50300 55462
rect 50356 55460 50380 55462
rect 50436 55460 50460 55462
rect 50516 55460 50540 55462
rect 50596 55460 50602 55462
rect 50294 55440 50602 55460
rect 50294 54428 50602 54448
rect 50294 54426 50300 54428
rect 50356 54426 50380 54428
rect 50436 54426 50460 54428
rect 50516 54426 50540 54428
rect 50596 54426 50602 54428
rect 50356 54374 50358 54426
rect 50538 54374 50540 54426
rect 50294 54372 50300 54374
rect 50356 54372 50380 54374
rect 50436 54372 50460 54374
rect 50516 54372 50540 54374
rect 50596 54372 50602 54374
rect 50294 54352 50602 54372
rect 50294 53340 50602 53360
rect 50294 53338 50300 53340
rect 50356 53338 50380 53340
rect 50436 53338 50460 53340
rect 50516 53338 50540 53340
rect 50596 53338 50602 53340
rect 50356 53286 50358 53338
rect 50538 53286 50540 53338
rect 50294 53284 50300 53286
rect 50356 53284 50380 53286
rect 50436 53284 50460 53286
rect 50516 53284 50540 53286
rect 50596 53284 50602 53286
rect 50294 53264 50602 53284
rect 50294 52252 50602 52272
rect 50294 52250 50300 52252
rect 50356 52250 50380 52252
rect 50436 52250 50460 52252
rect 50516 52250 50540 52252
rect 50596 52250 50602 52252
rect 50356 52198 50358 52250
rect 50538 52198 50540 52250
rect 50294 52196 50300 52198
rect 50356 52196 50380 52198
rect 50436 52196 50460 52198
rect 50516 52196 50540 52198
rect 50596 52196 50602 52198
rect 50294 52176 50602 52196
rect 50294 51164 50602 51184
rect 50294 51162 50300 51164
rect 50356 51162 50380 51164
rect 50436 51162 50460 51164
rect 50516 51162 50540 51164
rect 50596 51162 50602 51164
rect 50356 51110 50358 51162
rect 50538 51110 50540 51162
rect 50294 51108 50300 51110
rect 50356 51108 50380 51110
rect 50436 51108 50460 51110
rect 50516 51108 50540 51110
rect 50596 51108 50602 51110
rect 50294 51088 50602 51108
rect 50294 50076 50602 50096
rect 50294 50074 50300 50076
rect 50356 50074 50380 50076
rect 50436 50074 50460 50076
rect 50516 50074 50540 50076
rect 50596 50074 50602 50076
rect 50356 50022 50358 50074
rect 50538 50022 50540 50074
rect 50294 50020 50300 50022
rect 50356 50020 50380 50022
rect 50436 50020 50460 50022
rect 50516 50020 50540 50022
rect 50596 50020 50602 50022
rect 50294 50000 50602 50020
rect 50294 48988 50602 49008
rect 50294 48986 50300 48988
rect 50356 48986 50380 48988
rect 50436 48986 50460 48988
rect 50516 48986 50540 48988
rect 50596 48986 50602 48988
rect 50356 48934 50358 48986
rect 50538 48934 50540 48986
rect 50294 48932 50300 48934
rect 50356 48932 50380 48934
rect 50436 48932 50460 48934
rect 50516 48932 50540 48934
rect 50596 48932 50602 48934
rect 50294 48912 50602 48932
rect 50294 47900 50602 47920
rect 50294 47898 50300 47900
rect 50356 47898 50380 47900
rect 50436 47898 50460 47900
rect 50516 47898 50540 47900
rect 50596 47898 50602 47900
rect 50356 47846 50358 47898
rect 50538 47846 50540 47898
rect 50294 47844 50300 47846
rect 50356 47844 50380 47846
rect 50436 47844 50460 47846
rect 50516 47844 50540 47846
rect 50596 47844 50602 47846
rect 50294 47824 50602 47844
rect 50294 46812 50602 46832
rect 50294 46810 50300 46812
rect 50356 46810 50380 46812
rect 50436 46810 50460 46812
rect 50516 46810 50540 46812
rect 50596 46810 50602 46812
rect 50356 46758 50358 46810
rect 50538 46758 50540 46810
rect 50294 46756 50300 46758
rect 50356 46756 50380 46758
rect 50436 46756 50460 46758
rect 50516 46756 50540 46758
rect 50596 46756 50602 46758
rect 50294 46736 50602 46756
rect 50294 45724 50602 45744
rect 50294 45722 50300 45724
rect 50356 45722 50380 45724
rect 50436 45722 50460 45724
rect 50516 45722 50540 45724
rect 50596 45722 50602 45724
rect 50356 45670 50358 45722
rect 50538 45670 50540 45722
rect 50294 45668 50300 45670
rect 50356 45668 50380 45670
rect 50436 45668 50460 45670
rect 50516 45668 50540 45670
rect 50596 45668 50602 45670
rect 50294 45648 50602 45668
rect 50294 44636 50602 44656
rect 50294 44634 50300 44636
rect 50356 44634 50380 44636
rect 50436 44634 50460 44636
rect 50516 44634 50540 44636
rect 50596 44634 50602 44636
rect 50356 44582 50358 44634
rect 50538 44582 50540 44634
rect 50294 44580 50300 44582
rect 50356 44580 50380 44582
rect 50436 44580 50460 44582
rect 50516 44580 50540 44582
rect 50596 44580 50602 44582
rect 50294 44560 50602 44580
rect 50294 43548 50602 43568
rect 50294 43546 50300 43548
rect 50356 43546 50380 43548
rect 50436 43546 50460 43548
rect 50516 43546 50540 43548
rect 50596 43546 50602 43548
rect 50356 43494 50358 43546
rect 50538 43494 50540 43546
rect 50294 43492 50300 43494
rect 50356 43492 50380 43494
rect 50436 43492 50460 43494
rect 50516 43492 50540 43494
rect 50596 43492 50602 43494
rect 50294 43472 50602 43492
rect 50294 42460 50602 42480
rect 50294 42458 50300 42460
rect 50356 42458 50380 42460
rect 50436 42458 50460 42460
rect 50516 42458 50540 42460
rect 50596 42458 50602 42460
rect 50356 42406 50358 42458
rect 50538 42406 50540 42458
rect 50294 42404 50300 42406
rect 50356 42404 50380 42406
rect 50436 42404 50460 42406
rect 50516 42404 50540 42406
rect 50596 42404 50602 42406
rect 50294 42384 50602 42404
rect 50294 41372 50602 41392
rect 50294 41370 50300 41372
rect 50356 41370 50380 41372
rect 50436 41370 50460 41372
rect 50516 41370 50540 41372
rect 50596 41370 50602 41372
rect 50356 41318 50358 41370
rect 50538 41318 50540 41370
rect 50294 41316 50300 41318
rect 50356 41316 50380 41318
rect 50436 41316 50460 41318
rect 50516 41316 50540 41318
rect 50596 41316 50602 41318
rect 50294 41296 50602 41316
rect 50294 40284 50602 40304
rect 50294 40282 50300 40284
rect 50356 40282 50380 40284
rect 50436 40282 50460 40284
rect 50516 40282 50540 40284
rect 50596 40282 50602 40284
rect 50356 40230 50358 40282
rect 50538 40230 50540 40282
rect 50294 40228 50300 40230
rect 50356 40228 50380 40230
rect 50436 40228 50460 40230
rect 50516 40228 50540 40230
rect 50596 40228 50602 40230
rect 50294 40208 50602 40228
rect 50294 39196 50602 39216
rect 50294 39194 50300 39196
rect 50356 39194 50380 39196
rect 50436 39194 50460 39196
rect 50516 39194 50540 39196
rect 50596 39194 50602 39196
rect 50356 39142 50358 39194
rect 50538 39142 50540 39194
rect 50294 39140 50300 39142
rect 50356 39140 50380 39142
rect 50436 39140 50460 39142
rect 50516 39140 50540 39142
rect 50596 39140 50602 39142
rect 50294 39120 50602 39140
rect 50294 38108 50602 38128
rect 50294 38106 50300 38108
rect 50356 38106 50380 38108
rect 50436 38106 50460 38108
rect 50516 38106 50540 38108
rect 50596 38106 50602 38108
rect 50356 38054 50358 38106
rect 50538 38054 50540 38106
rect 50294 38052 50300 38054
rect 50356 38052 50380 38054
rect 50436 38052 50460 38054
rect 50516 38052 50540 38054
rect 50596 38052 50602 38054
rect 50294 38032 50602 38052
rect 50294 37020 50602 37040
rect 50294 37018 50300 37020
rect 50356 37018 50380 37020
rect 50436 37018 50460 37020
rect 50516 37018 50540 37020
rect 50596 37018 50602 37020
rect 50356 36966 50358 37018
rect 50538 36966 50540 37018
rect 50294 36964 50300 36966
rect 50356 36964 50380 36966
rect 50436 36964 50460 36966
rect 50516 36964 50540 36966
rect 50596 36964 50602 36966
rect 50294 36944 50602 36964
rect 50294 35932 50602 35952
rect 50294 35930 50300 35932
rect 50356 35930 50380 35932
rect 50436 35930 50460 35932
rect 50516 35930 50540 35932
rect 50596 35930 50602 35932
rect 50356 35878 50358 35930
rect 50538 35878 50540 35930
rect 50294 35876 50300 35878
rect 50356 35876 50380 35878
rect 50436 35876 50460 35878
rect 50516 35876 50540 35878
rect 50596 35876 50602 35878
rect 50294 35856 50602 35876
rect 50294 34844 50602 34864
rect 50294 34842 50300 34844
rect 50356 34842 50380 34844
rect 50436 34842 50460 34844
rect 50516 34842 50540 34844
rect 50596 34842 50602 34844
rect 50356 34790 50358 34842
rect 50538 34790 50540 34842
rect 50294 34788 50300 34790
rect 50356 34788 50380 34790
rect 50436 34788 50460 34790
rect 50516 34788 50540 34790
rect 50596 34788 50602 34790
rect 50294 34768 50602 34788
rect 50294 33756 50602 33776
rect 50294 33754 50300 33756
rect 50356 33754 50380 33756
rect 50436 33754 50460 33756
rect 50516 33754 50540 33756
rect 50596 33754 50602 33756
rect 50356 33702 50358 33754
rect 50538 33702 50540 33754
rect 50294 33700 50300 33702
rect 50356 33700 50380 33702
rect 50436 33700 50460 33702
rect 50516 33700 50540 33702
rect 50596 33700 50602 33702
rect 50294 33680 50602 33700
rect 50294 32668 50602 32688
rect 50294 32666 50300 32668
rect 50356 32666 50380 32668
rect 50436 32666 50460 32668
rect 50516 32666 50540 32668
rect 50596 32666 50602 32668
rect 50356 32614 50358 32666
rect 50538 32614 50540 32666
rect 50294 32612 50300 32614
rect 50356 32612 50380 32614
rect 50436 32612 50460 32614
rect 50516 32612 50540 32614
rect 50596 32612 50602 32614
rect 50294 32592 50602 32612
rect 50294 31580 50602 31600
rect 50294 31578 50300 31580
rect 50356 31578 50380 31580
rect 50436 31578 50460 31580
rect 50516 31578 50540 31580
rect 50596 31578 50602 31580
rect 50356 31526 50358 31578
rect 50538 31526 50540 31578
rect 50294 31524 50300 31526
rect 50356 31524 50380 31526
rect 50436 31524 50460 31526
rect 50516 31524 50540 31526
rect 50596 31524 50602 31526
rect 50294 31504 50602 31524
rect 50294 30492 50602 30512
rect 50294 30490 50300 30492
rect 50356 30490 50380 30492
rect 50436 30490 50460 30492
rect 50516 30490 50540 30492
rect 50596 30490 50602 30492
rect 50356 30438 50358 30490
rect 50538 30438 50540 30490
rect 50294 30436 50300 30438
rect 50356 30436 50380 30438
rect 50436 30436 50460 30438
rect 50516 30436 50540 30438
rect 50596 30436 50602 30438
rect 50294 30416 50602 30436
rect 50294 29404 50602 29424
rect 50294 29402 50300 29404
rect 50356 29402 50380 29404
rect 50436 29402 50460 29404
rect 50516 29402 50540 29404
rect 50596 29402 50602 29404
rect 50356 29350 50358 29402
rect 50538 29350 50540 29402
rect 50294 29348 50300 29350
rect 50356 29348 50380 29350
rect 50436 29348 50460 29350
rect 50516 29348 50540 29350
rect 50596 29348 50602 29350
rect 50294 29328 50602 29348
rect 50294 28316 50602 28336
rect 50294 28314 50300 28316
rect 50356 28314 50380 28316
rect 50436 28314 50460 28316
rect 50516 28314 50540 28316
rect 50596 28314 50602 28316
rect 50356 28262 50358 28314
rect 50538 28262 50540 28314
rect 50294 28260 50300 28262
rect 50356 28260 50380 28262
rect 50436 28260 50460 28262
rect 50516 28260 50540 28262
rect 50596 28260 50602 28262
rect 50294 28240 50602 28260
rect 50294 27228 50602 27248
rect 50294 27226 50300 27228
rect 50356 27226 50380 27228
rect 50436 27226 50460 27228
rect 50516 27226 50540 27228
rect 50596 27226 50602 27228
rect 50356 27174 50358 27226
rect 50538 27174 50540 27226
rect 50294 27172 50300 27174
rect 50356 27172 50380 27174
rect 50436 27172 50460 27174
rect 50516 27172 50540 27174
rect 50596 27172 50602 27174
rect 50294 27152 50602 27172
rect 50294 26140 50602 26160
rect 50294 26138 50300 26140
rect 50356 26138 50380 26140
rect 50436 26138 50460 26140
rect 50516 26138 50540 26140
rect 50596 26138 50602 26140
rect 50356 26086 50358 26138
rect 50538 26086 50540 26138
rect 50294 26084 50300 26086
rect 50356 26084 50380 26086
rect 50436 26084 50460 26086
rect 50516 26084 50540 26086
rect 50596 26084 50602 26086
rect 50294 26064 50602 26084
rect 50294 25052 50602 25072
rect 50294 25050 50300 25052
rect 50356 25050 50380 25052
rect 50436 25050 50460 25052
rect 50516 25050 50540 25052
rect 50596 25050 50602 25052
rect 50356 24998 50358 25050
rect 50538 24998 50540 25050
rect 50294 24996 50300 24998
rect 50356 24996 50380 24998
rect 50436 24996 50460 24998
rect 50516 24996 50540 24998
rect 50596 24996 50602 24998
rect 50294 24976 50602 24996
rect 50294 23964 50602 23984
rect 50294 23962 50300 23964
rect 50356 23962 50380 23964
rect 50436 23962 50460 23964
rect 50516 23962 50540 23964
rect 50596 23962 50602 23964
rect 50356 23910 50358 23962
rect 50538 23910 50540 23962
rect 50294 23908 50300 23910
rect 50356 23908 50380 23910
rect 50436 23908 50460 23910
rect 50516 23908 50540 23910
rect 50596 23908 50602 23910
rect 50294 23888 50602 23908
rect 50294 22876 50602 22896
rect 50294 22874 50300 22876
rect 50356 22874 50380 22876
rect 50436 22874 50460 22876
rect 50516 22874 50540 22876
rect 50596 22874 50602 22876
rect 50356 22822 50358 22874
rect 50538 22822 50540 22874
rect 50294 22820 50300 22822
rect 50356 22820 50380 22822
rect 50436 22820 50460 22822
rect 50516 22820 50540 22822
rect 50596 22820 50602 22822
rect 50294 22800 50602 22820
rect 50294 21788 50602 21808
rect 50294 21786 50300 21788
rect 50356 21786 50380 21788
rect 50436 21786 50460 21788
rect 50516 21786 50540 21788
rect 50596 21786 50602 21788
rect 50356 21734 50358 21786
rect 50538 21734 50540 21786
rect 50294 21732 50300 21734
rect 50356 21732 50380 21734
rect 50436 21732 50460 21734
rect 50516 21732 50540 21734
rect 50596 21732 50602 21734
rect 50294 21712 50602 21732
rect 50294 20700 50602 20720
rect 50294 20698 50300 20700
rect 50356 20698 50380 20700
rect 50436 20698 50460 20700
rect 50516 20698 50540 20700
rect 50596 20698 50602 20700
rect 50356 20646 50358 20698
rect 50538 20646 50540 20698
rect 50294 20644 50300 20646
rect 50356 20644 50380 20646
rect 50436 20644 50460 20646
rect 50516 20644 50540 20646
rect 50596 20644 50602 20646
rect 50294 20624 50602 20644
rect 50294 19612 50602 19632
rect 50294 19610 50300 19612
rect 50356 19610 50380 19612
rect 50436 19610 50460 19612
rect 50516 19610 50540 19612
rect 50596 19610 50602 19612
rect 50356 19558 50358 19610
rect 50538 19558 50540 19610
rect 50294 19556 50300 19558
rect 50356 19556 50380 19558
rect 50436 19556 50460 19558
rect 50516 19556 50540 19558
rect 50596 19556 50602 19558
rect 50294 19536 50602 19556
rect 50294 18524 50602 18544
rect 50294 18522 50300 18524
rect 50356 18522 50380 18524
rect 50436 18522 50460 18524
rect 50516 18522 50540 18524
rect 50596 18522 50602 18524
rect 50356 18470 50358 18522
rect 50538 18470 50540 18522
rect 50294 18468 50300 18470
rect 50356 18468 50380 18470
rect 50436 18468 50460 18470
rect 50516 18468 50540 18470
rect 50596 18468 50602 18470
rect 50294 18448 50602 18468
rect 50294 17436 50602 17456
rect 50294 17434 50300 17436
rect 50356 17434 50380 17436
rect 50436 17434 50460 17436
rect 50516 17434 50540 17436
rect 50596 17434 50602 17436
rect 50356 17382 50358 17434
rect 50538 17382 50540 17434
rect 50294 17380 50300 17382
rect 50356 17380 50380 17382
rect 50436 17380 50460 17382
rect 50516 17380 50540 17382
rect 50596 17380 50602 17382
rect 50294 17360 50602 17380
rect 63052 16590 63080 59910
rect 63880 58954 63908 117234
rect 64064 117094 64092 119326
rect 66994 119326 67312 119354
rect 66994 119200 67050 119326
rect 67284 117162 67312 119326
rect 70858 119200 70914 120000
rect 74722 119354 74778 120000
rect 74722 119326 75040 119354
rect 74722 119200 74778 119326
rect 70872 117298 70900 119200
rect 70860 117292 70912 117298
rect 70860 117234 70912 117240
rect 75012 117162 75040 119326
rect 78586 119200 78642 120000
rect 77206 118416 77262 118425
rect 77206 118351 77262 118360
rect 66536 117156 66588 117162
rect 66536 117098 66588 117104
rect 67272 117156 67324 117162
rect 67272 117098 67324 117104
rect 75000 117156 75052 117162
rect 75000 117098 75052 117104
rect 64052 117088 64104 117094
rect 64052 117030 64104 117036
rect 65654 116988 65962 117008
rect 65654 116986 65660 116988
rect 65716 116986 65740 116988
rect 65796 116986 65820 116988
rect 65876 116986 65900 116988
rect 65956 116986 65962 116988
rect 65716 116934 65718 116986
rect 65898 116934 65900 116986
rect 65654 116932 65660 116934
rect 65716 116932 65740 116934
rect 65796 116932 65820 116934
rect 65876 116932 65900 116934
rect 65956 116932 65962 116934
rect 65654 116912 65962 116932
rect 65654 115900 65962 115920
rect 65654 115898 65660 115900
rect 65716 115898 65740 115900
rect 65796 115898 65820 115900
rect 65876 115898 65900 115900
rect 65956 115898 65962 115900
rect 65716 115846 65718 115898
rect 65898 115846 65900 115898
rect 65654 115844 65660 115846
rect 65716 115844 65740 115846
rect 65796 115844 65820 115846
rect 65876 115844 65900 115846
rect 65956 115844 65962 115846
rect 65654 115824 65962 115844
rect 65654 114812 65962 114832
rect 65654 114810 65660 114812
rect 65716 114810 65740 114812
rect 65796 114810 65820 114812
rect 65876 114810 65900 114812
rect 65956 114810 65962 114812
rect 65716 114758 65718 114810
rect 65898 114758 65900 114810
rect 65654 114756 65660 114758
rect 65716 114756 65740 114758
rect 65796 114756 65820 114758
rect 65876 114756 65900 114758
rect 65956 114756 65962 114758
rect 65654 114736 65962 114756
rect 65654 113724 65962 113744
rect 65654 113722 65660 113724
rect 65716 113722 65740 113724
rect 65796 113722 65820 113724
rect 65876 113722 65900 113724
rect 65956 113722 65962 113724
rect 65716 113670 65718 113722
rect 65898 113670 65900 113722
rect 65654 113668 65660 113670
rect 65716 113668 65740 113670
rect 65796 113668 65820 113670
rect 65876 113668 65900 113670
rect 65956 113668 65962 113670
rect 65654 113648 65962 113668
rect 65654 112636 65962 112656
rect 65654 112634 65660 112636
rect 65716 112634 65740 112636
rect 65796 112634 65820 112636
rect 65876 112634 65900 112636
rect 65956 112634 65962 112636
rect 65716 112582 65718 112634
rect 65898 112582 65900 112634
rect 65654 112580 65660 112582
rect 65716 112580 65740 112582
rect 65796 112580 65820 112582
rect 65876 112580 65900 112582
rect 65956 112580 65962 112582
rect 65654 112560 65962 112580
rect 66548 111926 66576 117098
rect 66720 117088 66772 117094
rect 66720 117030 66772 117036
rect 71320 117088 71372 117094
rect 71320 117030 71372 117036
rect 74540 117088 74592 117094
rect 74540 117030 74592 117036
rect 66732 116890 66760 117030
rect 66720 116884 66772 116890
rect 66720 116826 66772 116832
rect 66536 111920 66588 111926
rect 66536 111862 66588 111868
rect 65654 111548 65962 111568
rect 65654 111546 65660 111548
rect 65716 111546 65740 111548
rect 65796 111546 65820 111548
rect 65876 111546 65900 111548
rect 65956 111546 65962 111548
rect 65716 111494 65718 111546
rect 65898 111494 65900 111546
rect 65654 111492 65660 111494
rect 65716 111492 65740 111494
rect 65796 111492 65820 111494
rect 65876 111492 65900 111494
rect 65956 111492 65962 111494
rect 65654 111472 65962 111492
rect 65654 110460 65962 110480
rect 65654 110458 65660 110460
rect 65716 110458 65740 110460
rect 65796 110458 65820 110460
rect 65876 110458 65900 110460
rect 65956 110458 65962 110460
rect 65716 110406 65718 110458
rect 65898 110406 65900 110458
rect 65654 110404 65660 110406
rect 65716 110404 65740 110406
rect 65796 110404 65820 110406
rect 65876 110404 65900 110406
rect 65956 110404 65962 110406
rect 65654 110384 65962 110404
rect 65654 109372 65962 109392
rect 65654 109370 65660 109372
rect 65716 109370 65740 109372
rect 65796 109370 65820 109372
rect 65876 109370 65900 109372
rect 65956 109370 65962 109372
rect 65716 109318 65718 109370
rect 65898 109318 65900 109370
rect 65654 109316 65660 109318
rect 65716 109316 65740 109318
rect 65796 109316 65820 109318
rect 65876 109316 65900 109318
rect 65956 109316 65962 109318
rect 65654 109296 65962 109316
rect 65654 108284 65962 108304
rect 65654 108282 65660 108284
rect 65716 108282 65740 108284
rect 65796 108282 65820 108284
rect 65876 108282 65900 108284
rect 65956 108282 65962 108284
rect 65716 108230 65718 108282
rect 65898 108230 65900 108282
rect 65654 108228 65660 108230
rect 65716 108228 65740 108230
rect 65796 108228 65820 108230
rect 65876 108228 65900 108230
rect 65956 108228 65962 108230
rect 65654 108208 65962 108228
rect 65654 107196 65962 107216
rect 65654 107194 65660 107196
rect 65716 107194 65740 107196
rect 65796 107194 65820 107196
rect 65876 107194 65900 107196
rect 65956 107194 65962 107196
rect 65716 107142 65718 107194
rect 65898 107142 65900 107194
rect 65654 107140 65660 107142
rect 65716 107140 65740 107142
rect 65796 107140 65820 107142
rect 65876 107140 65900 107142
rect 65956 107140 65962 107142
rect 65654 107120 65962 107140
rect 65654 106108 65962 106128
rect 65654 106106 65660 106108
rect 65716 106106 65740 106108
rect 65796 106106 65820 106108
rect 65876 106106 65900 106108
rect 65956 106106 65962 106108
rect 65716 106054 65718 106106
rect 65898 106054 65900 106106
rect 65654 106052 65660 106054
rect 65716 106052 65740 106054
rect 65796 106052 65820 106054
rect 65876 106052 65900 106054
rect 65956 106052 65962 106054
rect 65654 106032 65962 106052
rect 65654 105020 65962 105040
rect 65654 105018 65660 105020
rect 65716 105018 65740 105020
rect 65796 105018 65820 105020
rect 65876 105018 65900 105020
rect 65956 105018 65962 105020
rect 65716 104966 65718 105018
rect 65898 104966 65900 105018
rect 65654 104964 65660 104966
rect 65716 104964 65740 104966
rect 65796 104964 65820 104966
rect 65876 104964 65900 104966
rect 65956 104964 65962 104966
rect 65654 104944 65962 104964
rect 65654 103932 65962 103952
rect 65654 103930 65660 103932
rect 65716 103930 65740 103932
rect 65796 103930 65820 103932
rect 65876 103930 65900 103932
rect 65956 103930 65962 103932
rect 65716 103878 65718 103930
rect 65898 103878 65900 103930
rect 65654 103876 65660 103878
rect 65716 103876 65740 103878
rect 65796 103876 65820 103878
rect 65876 103876 65900 103878
rect 65956 103876 65962 103878
rect 65654 103856 65962 103876
rect 65654 102844 65962 102864
rect 65654 102842 65660 102844
rect 65716 102842 65740 102844
rect 65796 102842 65820 102844
rect 65876 102842 65900 102844
rect 65956 102842 65962 102844
rect 65716 102790 65718 102842
rect 65898 102790 65900 102842
rect 65654 102788 65660 102790
rect 65716 102788 65740 102790
rect 65796 102788 65820 102790
rect 65876 102788 65900 102790
rect 65956 102788 65962 102790
rect 65654 102768 65962 102788
rect 65654 101756 65962 101776
rect 65654 101754 65660 101756
rect 65716 101754 65740 101756
rect 65796 101754 65820 101756
rect 65876 101754 65900 101756
rect 65956 101754 65962 101756
rect 65716 101702 65718 101754
rect 65898 101702 65900 101754
rect 65654 101700 65660 101702
rect 65716 101700 65740 101702
rect 65796 101700 65820 101702
rect 65876 101700 65900 101702
rect 65956 101700 65962 101702
rect 65654 101680 65962 101700
rect 65654 100668 65962 100688
rect 65654 100666 65660 100668
rect 65716 100666 65740 100668
rect 65796 100666 65820 100668
rect 65876 100666 65900 100668
rect 65956 100666 65962 100668
rect 65716 100614 65718 100666
rect 65898 100614 65900 100666
rect 65654 100612 65660 100614
rect 65716 100612 65740 100614
rect 65796 100612 65820 100614
rect 65876 100612 65900 100614
rect 65956 100612 65962 100614
rect 65654 100592 65962 100612
rect 65654 99580 65962 99600
rect 65654 99578 65660 99580
rect 65716 99578 65740 99580
rect 65796 99578 65820 99580
rect 65876 99578 65900 99580
rect 65956 99578 65962 99580
rect 65716 99526 65718 99578
rect 65898 99526 65900 99578
rect 65654 99524 65660 99526
rect 65716 99524 65740 99526
rect 65796 99524 65820 99526
rect 65876 99524 65900 99526
rect 65956 99524 65962 99526
rect 65654 99504 65962 99524
rect 65654 98492 65962 98512
rect 65654 98490 65660 98492
rect 65716 98490 65740 98492
rect 65796 98490 65820 98492
rect 65876 98490 65900 98492
rect 65956 98490 65962 98492
rect 65716 98438 65718 98490
rect 65898 98438 65900 98490
rect 65654 98436 65660 98438
rect 65716 98436 65740 98438
rect 65796 98436 65820 98438
rect 65876 98436 65900 98438
rect 65956 98436 65962 98438
rect 65654 98416 65962 98436
rect 65654 97404 65962 97424
rect 65654 97402 65660 97404
rect 65716 97402 65740 97404
rect 65796 97402 65820 97404
rect 65876 97402 65900 97404
rect 65956 97402 65962 97404
rect 65716 97350 65718 97402
rect 65898 97350 65900 97402
rect 65654 97348 65660 97350
rect 65716 97348 65740 97350
rect 65796 97348 65820 97350
rect 65876 97348 65900 97350
rect 65956 97348 65962 97350
rect 65654 97328 65962 97348
rect 65654 96316 65962 96336
rect 65654 96314 65660 96316
rect 65716 96314 65740 96316
rect 65796 96314 65820 96316
rect 65876 96314 65900 96316
rect 65956 96314 65962 96316
rect 65716 96262 65718 96314
rect 65898 96262 65900 96314
rect 65654 96260 65660 96262
rect 65716 96260 65740 96262
rect 65796 96260 65820 96262
rect 65876 96260 65900 96262
rect 65956 96260 65962 96262
rect 65654 96240 65962 96260
rect 65654 95228 65962 95248
rect 65654 95226 65660 95228
rect 65716 95226 65740 95228
rect 65796 95226 65820 95228
rect 65876 95226 65900 95228
rect 65956 95226 65962 95228
rect 65716 95174 65718 95226
rect 65898 95174 65900 95226
rect 65654 95172 65660 95174
rect 65716 95172 65740 95174
rect 65796 95172 65820 95174
rect 65876 95172 65900 95174
rect 65956 95172 65962 95174
rect 65654 95152 65962 95172
rect 65654 94140 65962 94160
rect 65654 94138 65660 94140
rect 65716 94138 65740 94140
rect 65796 94138 65820 94140
rect 65876 94138 65900 94140
rect 65956 94138 65962 94140
rect 65716 94086 65718 94138
rect 65898 94086 65900 94138
rect 65654 94084 65660 94086
rect 65716 94084 65740 94086
rect 65796 94084 65820 94086
rect 65876 94084 65900 94086
rect 65956 94084 65962 94086
rect 65654 94064 65962 94084
rect 65654 93052 65962 93072
rect 65654 93050 65660 93052
rect 65716 93050 65740 93052
rect 65796 93050 65820 93052
rect 65876 93050 65900 93052
rect 65956 93050 65962 93052
rect 65716 92998 65718 93050
rect 65898 92998 65900 93050
rect 65654 92996 65660 92998
rect 65716 92996 65740 92998
rect 65796 92996 65820 92998
rect 65876 92996 65900 92998
rect 65956 92996 65962 92998
rect 65654 92976 65962 92996
rect 65654 91964 65962 91984
rect 65654 91962 65660 91964
rect 65716 91962 65740 91964
rect 65796 91962 65820 91964
rect 65876 91962 65900 91964
rect 65956 91962 65962 91964
rect 65716 91910 65718 91962
rect 65898 91910 65900 91962
rect 65654 91908 65660 91910
rect 65716 91908 65740 91910
rect 65796 91908 65820 91910
rect 65876 91908 65900 91910
rect 65956 91908 65962 91910
rect 65654 91888 65962 91908
rect 65654 90876 65962 90896
rect 65654 90874 65660 90876
rect 65716 90874 65740 90876
rect 65796 90874 65820 90876
rect 65876 90874 65900 90876
rect 65956 90874 65962 90876
rect 65716 90822 65718 90874
rect 65898 90822 65900 90874
rect 65654 90820 65660 90822
rect 65716 90820 65740 90822
rect 65796 90820 65820 90822
rect 65876 90820 65900 90822
rect 65956 90820 65962 90822
rect 65654 90800 65962 90820
rect 65654 89788 65962 89808
rect 65654 89786 65660 89788
rect 65716 89786 65740 89788
rect 65796 89786 65820 89788
rect 65876 89786 65900 89788
rect 65956 89786 65962 89788
rect 65716 89734 65718 89786
rect 65898 89734 65900 89786
rect 65654 89732 65660 89734
rect 65716 89732 65740 89734
rect 65796 89732 65820 89734
rect 65876 89732 65900 89734
rect 65956 89732 65962 89734
rect 65654 89712 65962 89732
rect 65654 88700 65962 88720
rect 65654 88698 65660 88700
rect 65716 88698 65740 88700
rect 65796 88698 65820 88700
rect 65876 88698 65900 88700
rect 65956 88698 65962 88700
rect 65716 88646 65718 88698
rect 65898 88646 65900 88698
rect 65654 88644 65660 88646
rect 65716 88644 65740 88646
rect 65796 88644 65820 88646
rect 65876 88644 65900 88646
rect 65956 88644 65962 88646
rect 65654 88624 65962 88644
rect 65654 87612 65962 87632
rect 65654 87610 65660 87612
rect 65716 87610 65740 87612
rect 65796 87610 65820 87612
rect 65876 87610 65900 87612
rect 65956 87610 65962 87612
rect 65716 87558 65718 87610
rect 65898 87558 65900 87610
rect 65654 87556 65660 87558
rect 65716 87556 65740 87558
rect 65796 87556 65820 87558
rect 65876 87556 65900 87558
rect 65956 87556 65962 87558
rect 65654 87536 65962 87556
rect 65654 86524 65962 86544
rect 65654 86522 65660 86524
rect 65716 86522 65740 86524
rect 65796 86522 65820 86524
rect 65876 86522 65900 86524
rect 65956 86522 65962 86524
rect 65716 86470 65718 86522
rect 65898 86470 65900 86522
rect 65654 86468 65660 86470
rect 65716 86468 65740 86470
rect 65796 86468 65820 86470
rect 65876 86468 65900 86470
rect 65956 86468 65962 86470
rect 65654 86448 65962 86468
rect 65654 85436 65962 85456
rect 65654 85434 65660 85436
rect 65716 85434 65740 85436
rect 65796 85434 65820 85436
rect 65876 85434 65900 85436
rect 65956 85434 65962 85436
rect 65716 85382 65718 85434
rect 65898 85382 65900 85434
rect 65654 85380 65660 85382
rect 65716 85380 65740 85382
rect 65796 85380 65820 85382
rect 65876 85380 65900 85382
rect 65956 85380 65962 85382
rect 65654 85360 65962 85380
rect 65654 84348 65962 84368
rect 65654 84346 65660 84348
rect 65716 84346 65740 84348
rect 65796 84346 65820 84348
rect 65876 84346 65900 84348
rect 65956 84346 65962 84348
rect 65716 84294 65718 84346
rect 65898 84294 65900 84346
rect 65654 84292 65660 84294
rect 65716 84292 65740 84294
rect 65796 84292 65820 84294
rect 65876 84292 65900 84294
rect 65956 84292 65962 84294
rect 65654 84272 65962 84292
rect 65654 83260 65962 83280
rect 65654 83258 65660 83260
rect 65716 83258 65740 83260
rect 65796 83258 65820 83260
rect 65876 83258 65900 83260
rect 65956 83258 65962 83260
rect 65716 83206 65718 83258
rect 65898 83206 65900 83258
rect 65654 83204 65660 83206
rect 65716 83204 65740 83206
rect 65796 83204 65820 83206
rect 65876 83204 65900 83206
rect 65956 83204 65962 83206
rect 65654 83184 65962 83204
rect 65654 82172 65962 82192
rect 65654 82170 65660 82172
rect 65716 82170 65740 82172
rect 65796 82170 65820 82172
rect 65876 82170 65900 82172
rect 65956 82170 65962 82172
rect 65716 82118 65718 82170
rect 65898 82118 65900 82170
rect 65654 82116 65660 82118
rect 65716 82116 65740 82118
rect 65796 82116 65820 82118
rect 65876 82116 65900 82118
rect 65956 82116 65962 82118
rect 65654 82096 65962 82116
rect 65654 81084 65962 81104
rect 65654 81082 65660 81084
rect 65716 81082 65740 81084
rect 65796 81082 65820 81084
rect 65876 81082 65900 81084
rect 65956 81082 65962 81084
rect 65716 81030 65718 81082
rect 65898 81030 65900 81082
rect 65654 81028 65660 81030
rect 65716 81028 65740 81030
rect 65796 81028 65820 81030
rect 65876 81028 65900 81030
rect 65956 81028 65962 81030
rect 65654 81008 65962 81028
rect 65654 79996 65962 80016
rect 65654 79994 65660 79996
rect 65716 79994 65740 79996
rect 65796 79994 65820 79996
rect 65876 79994 65900 79996
rect 65956 79994 65962 79996
rect 65716 79942 65718 79994
rect 65898 79942 65900 79994
rect 65654 79940 65660 79942
rect 65716 79940 65740 79942
rect 65796 79940 65820 79942
rect 65876 79940 65900 79942
rect 65956 79940 65962 79942
rect 65654 79920 65962 79940
rect 65654 78908 65962 78928
rect 65654 78906 65660 78908
rect 65716 78906 65740 78908
rect 65796 78906 65820 78908
rect 65876 78906 65900 78908
rect 65956 78906 65962 78908
rect 65716 78854 65718 78906
rect 65898 78854 65900 78906
rect 65654 78852 65660 78854
rect 65716 78852 65740 78854
rect 65796 78852 65820 78854
rect 65876 78852 65900 78854
rect 65956 78852 65962 78854
rect 65654 78832 65962 78852
rect 65654 77820 65962 77840
rect 65654 77818 65660 77820
rect 65716 77818 65740 77820
rect 65796 77818 65820 77820
rect 65876 77818 65900 77820
rect 65956 77818 65962 77820
rect 65716 77766 65718 77818
rect 65898 77766 65900 77818
rect 65654 77764 65660 77766
rect 65716 77764 65740 77766
rect 65796 77764 65820 77766
rect 65876 77764 65900 77766
rect 65956 77764 65962 77766
rect 65654 77744 65962 77764
rect 65654 76732 65962 76752
rect 65654 76730 65660 76732
rect 65716 76730 65740 76732
rect 65796 76730 65820 76732
rect 65876 76730 65900 76732
rect 65956 76730 65962 76732
rect 65716 76678 65718 76730
rect 65898 76678 65900 76730
rect 65654 76676 65660 76678
rect 65716 76676 65740 76678
rect 65796 76676 65820 76678
rect 65876 76676 65900 76678
rect 65956 76676 65962 76678
rect 65654 76656 65962 76676
rect 65654 75644 65962 75664
rect 65654 75642 65660 75644
rect 65716 75642 65740 75644
rect 65796 75642 65820 75644
rect 65876 75642 65900 75644
rect 65956 75642 65962 75644
rect 65716 75590 65718 75642
rect 65898 75590 65900 75642
rect 65654 75588 65660 75590
rect 65716 75588 65740 75590
rect 65796 75588 65820 75590
rect 65876 75588 65900 75590
rect 65956 75588 65962 75590
rect 65654 75568 65962 75588
rect 65654 74556 65962 74576
rect 65654 74554 65660 74556
rect 65716 74554 65740 74556
rect 65796 74554 65820 74556
rect 65876 74554 65900 74556
rect 65956 74554 65962 74556
rect 65716 74502 65718 74554
rect 65898 74502 65900 74554
rect 65654 74500 65660 74502
rect 65716 74500 65740 74502
rect 65796 74500 65820 74502
rect 65876 74500 65900 74502
rect 65956 74500 65962 74502
rect 65654 74480 65962 74500
rect 65654 73468 65962 73488
rect 65654 73466 65660 73468
rect 65716 73466 65740 73468
rect 65796 73466 65820 73468
rect 65876 73466 65900 73468
rect 65956 73466 65962 73468
rect 65716 73414 65718 73466
rect 65898 73414 65900 73466
rect 65654 73412 65660 73414
rect 65716 73412 65740 73414
rect 65796 73412 65820 73414
rect 65876 73412 65900 73414
rect 65956 73412 65962 73414
rect 65654 73392 65962 73412
rect 65654 72380 65962 72400
rect 65654 72378 65660 72380
rect 65716 72378 65740 72380
rect 65796 72378 65820 72380
rect 65876 72378 65900 72380
rect 65956 72378 65962 72380
rect 65716 72326 65718 72378
rect 65898 72326 65900 72378
rect 65654 72324 65660 72326
rect 65716 72324 65740 72326
rect 65796 72324 65820 72326
rect 65876 72324 65900 72326
rect 65956 72324 65962 72326
rect 65654 72304 65962 72324
rect 65654 71292 65962 71312
rect 65654 71290 65660 71292
rect 65716 71290 65740 71292
rect 65796 71290 65820 71292
rect 65876 71290 65900 71292
rect 65956 71290 65962 71292
rect 65716 71238 65718 71290
rect 65898 71238 65900 71290
rect 65654 71236 65660 71238
rect 65716 71236 65740 71238
rect 65796 71236 65820 71238
rect 65876 71236 65900 71238
rect 65956 71236 65962 71238
rect 65654 71216 65962 71236
rect 65654 70204 65962 70224
rect 65654 70202 65660 70204
rect 65716 70202 65740 70204
rect 65796 70202 65820 70204
rect 65876 70202 65900 70204
rect 65956 70202 65962 70204
rect 65716 70150 65718 70202
rect 65898 70150 65900 70202
rect 65654 70148 65660 70150
rect 65716 70148 65740 70150
rect 65796 70148 65820 70150
rect 65876 70148 65900 70150
rect 65956 70148 65962 70150
rect 65654 70128 65962 70148
rect 65654 69116 65962 69136
rect 65654 69114 65660 69116
rect 65716 69114 65740 69116
rect 65796 69114 65820 69116
rect 65876 69114 65900 69116
rect 65956 69114 65962 69116
rect 65716 69062 65718 69114
rect 65898 69062 65900 69114
rect 65654 69060 65660 69062
rect 65716 69060 65740 69062
rect 65796 69060 65820 69062
rect 65876 69060 65900 69062
rect 65956 69060 65962 69062
rect 65654 69040 65962 69060
rect 65654 68028 65962 68048
rect 65654 68026 65660 68028
rect 65716 68026 65740 68028
rect 65796 68026 65820 68028
rect 65876 68026 65900 68028
rect 65956 68026 65962 68028
rect 65716 67974 65718 68026
rect 65898 67974 65900 68026
rect 65654 67972 65660 67974
rect 65716 67972 65740 67974
rect 65796 67972 65820 67974
rect 65876 67972 65900 67974
rect 65956 67972 65962 67974
rect 65654 67952 65962 67972
rect 65654 66940 65962 66960
rect 65654 66938 65660 66940
rect 65716 66938 65740 66940
rect 65796 66938 65820 66940
rect 65876 66938 65900 66940
rect 65956 66938 65962 66940
rect 65716 66886 65718 66938
rect 65898 66886 65900 66938
rect 65654 66884 65660 66886
rect 65716 66884 65740 66886
rect 65796 66884 65820 66886
rect 65876 66884 65900 66886
rect 65956 66884 65962 66886
rect 65654 66864 65962 66884
rect 65654 65852 65962 65872
rect 65654 65850 65660 65852
rect 65716 65850 65740 65852
rect 65796 65850 65820 65852
rect 65876 65850 65900 65852
rect 65956 65850 65962 65852
rect 65716 65798 65718 65850
rect 65898 65798 65900 65850
rect 65654 65796 65660 65798
rect 65716 65796 65740 65798
rect 65796 65796 65820 65798
rect 65876 65796 65900 65798
rect 65956 65796 65962 65798
rect 65654 65776 65962 65796
rect 65654 64764 65962 64784
rect 65654 64762 65660 64764
rect 65716 64762 65740 64764
rect 65796 64762 65820 64764
rect 65876 64762 65900 64764
rect 65956 64762 65962 64764
rect 65716 64710 65718 64762
rect 65898 64710 65900 64762
rect 65654 64708 65660 64710
rect 65716 64708 65740 64710
rect 65796 64708 65820 64710
rect 65876 64708 65900 64710
rect 65956 64708 65962 64710
rect 65654 64688 65962 64708
rect 65654 63676 65962 63696
rect 65654 63674 65660 63676
rect 65716 63674 65740 63676
rect 65796 63674 65820 63676
rect 65876 63674 65900 63676
rect 65956 63674 65962 63676
rect 65716 63622 65718 63674
rect 65898 63622 65900 63674
rect 65654 63620 65660 63622
rect 65716 63620 65740 63622
rect 65796 63620 65820 63622
rect 65876 63620 65900 63622
rect 65956 63620 65962 63622
rect 65654 63600 65962 63620
rect 65654 62588 65962 62608
rect 65654 62586 65660 62588
rect 65716 62586 65740 62588
rect 65796 62586 65820 62588
rect 65876 62586 65900 62588
rect 65956 62586 65962 62588
rect 65716 62534 65718 62586
rect 65898 62534 65900 62586
rect 65654 62532 65660 62534
rect 65716 62532 65740 62534
rect 65796 62532 65820 62534
rect 65876 62532 65900 62534
rect 65956 62532 65962 62534
rect 65654 62512 65962 62532
rect 65654 61500 65962 61520
rect 65654 61498 65660 61500
rect 65716 61498 65740 61500
rect 65796 61498 65820 61500
rect 65876 61498 65900 61500
rect 65956 61498 65962 61500
rect 65716 61446 65718 61498
rect 65898 61446 65900 61498
rect 65654 61444 65660 61446
rect 65716 61444 65740 61446
rect 65796 61444 65820 61446
rect 65876 61444 65900 61446
rect 65956 61444 65962 61446
rect 65654 61424 65962 61444
rect 65654 60412 65962 60432
rect 65654 60410 65660 60412
rect 65716 60410 65740 60412
rect 65796 60410 65820 60412
rect 65876 60410 65900 60412
rect 65956 60410 65962 60412
rect 65716 60358 65718 60410
rect 65898 60358 65900 60410
rect 65654 60356 65660 60358
rect 65716 60356 65740 60358
rect 65796 60356 65820 60358
rect 65876 60356 65900 60358
rect 65956 60356 65962 60358
rect 65654 60336 65962 60356
rect 71332 59634 71360 117030
rect 74552 116754 74580 117030
rect 77220 116890 77248 118351
rect 78600 117298 78628 119200
rect 78588 117292 78640 117298
rect 78588 117234 78640 117240
rect 77944 117224 77996 117230
rect 77944 117166 77996 117172
rect 77208 116884 77260 116890
rect 77208 116826 77260 116832
rect 74540 116748 74592 116754
rect 74540 116690 74592 116696
rect 77852 116680 77904 116686
rect 77852 116622 77904 116628
rect 77864 116006 77892 116622
rect 77852 116000 77904 116006
rect 77852 115942 77904 115948
rect 77392 114504 77444 114510
rect 77392 114446 77444 114452
rect 76012 111852 76064 111858
rect 76012 111794 76064 111800
rect 76024 106418 76052 111794
rect 76012 106412 76064 106418
rect 76012 106354 76064 106360
rect 77300 103148 77352 103154
rect 77300 103090 77352 103096
rect 77312 102950 77340 103090
rect 77300 102944 77352 102950
rect 77300 102886 77352 102892
rect 76748 72072 76800 72078
rect 76748 72014 76800 72020
rect 76564 71596 76616 71602
rect 76564 71538 76616 71544
rect 76576 71194 76604 71538
rect 76564 71188 76616 71194
rect 76564 71130 76616 71136
rect 76760 70990 76788 72014
rect 76748 70984 76800 70990
rect 76748 70926 76800 70932
rect 77312 60654 77340 102886
rect 77300 60648 77352 60654
rect 77300 60590 77352 60596
rect 71320 59628 71372 59634
rect 71320 59570 71372 59576
rect 77404 59566 77432 114446
rect 77956 113174 77984 117166
rect 78036 114368 78088 114374
rect 78034 114336 78036 114345
rect 78088 114336 78090 114345
rect 78034 114271 78090 114280
rect 77956 113146 78076 113174
rect 77760 110764 77812 110770
rect 77760 110706 77812 110712
rect 77668 83564 77720 83570
rect 77668 83506 77720 83512
rect 77576 79212 77628 79218
rect 77576 79154 77628 79160
rect 77588 78985 77616 79154
rect 77574 78976 77630 78985
rect 77574 78911 77630 78920
rect 77680 74534 77708 83506
rect 77588 74506 77708 74534
rect 77484 69760 77536 69766
rect 77484 69702 77536 69708
rect 77496 59974 77524 69702
rect 77588 60518 77616 74506
rect 77668 70984 77720 70990
rect 77668 70926 77720 70932
rect 77576 60512 77628 60518
rect 77576 60454 77628 60460
rect 77484 59968 77536 59974
rect 77484 59910 77536 59916
rect 77392 59560 77444 59566
rect 77392 59502 77444 59508
rect 77392 59424 77444 59430
rect 77392 59366 77444 59372
rect 65654 59324 65962 59344
rect 65654 59322 65660 59324
rect 65716 59322 65740 59324
rect 65796 59322 65820 59324
rect 65876 59322 65900 59324
rect 65956 59322 65962 59324
rect 65716 59270 65718 59322
rect 65898 59270 65900 59322
rect 65654 59268 65660 59270
rect 65716 59268 65740 59270
rect 65796 59268 65820 59270
rect 65876 59268 65900 59270
rect 65956 59268 65962 59270
rect 65654 59248 65962 59268
rect 63868 58948 63920 58954
rect 63868 58890 63920 58896
rect 65654 58236 65962 58256
rect 65654 58234 65660 58236
rect 65716 58234 65740 58236
rect 65796 58234 65820 58236
rect 65876 58234 65900 58236
rect 65956 58234 65962 58236
rect 65716 58182 65718 58234
rect 65898 58182 65900 58234
rect 65654 58180 65660 58182
rect 65716 58180 65740 58182
rect 65796 58180 65820 58182
rect 65876 58180 65900 58182
rect 65956 58180 65962 58182
rect 65654 58160 65962 58180
rect 65654 57148 65962 57168
rect 65654 57146 65660 57148
rect 65716 57146 65740 57148
rect 65796 57146 65820 57148
rect 65876 57146 65900 57148
rect 65956 57146 65962 57148
rect 65716 57094 65718 57146
rect 65898 57094 65900 57146
rect 65654 57092 65660 57094
rect 65716 57092 65740 57094
rect 65796 57092 65820 57094
rect 65876 57092 65900 57094
rect 65956 57092 65962 57094
rect 65654 57072 65962 57092
rect 65654 56060 65962 56080
rect 65654 56058 65660 56060
rect 65716 56058 65740 56060
rect 65796 56058 65820 56060
rect 65876 56058 65900 56060
rect 65956 56058 65962 56060
rect 65716 56006 65718 56058
rect 65898 56006 65900 56058
rect 65654 56004 65660 56006
rect 65716 56004 65740 56006
rect 65796 56004 65820 56006
rect 65876 56004 65900 56006
rect 65956 56004 65962 56006
rect 65654 55984 65962 56004
rect 65654 54972 65962 54992
rect 65654 54970 65660 54972
rect 65716 54970 65740 54972
rect 65796 54970 65820 54972
rect 65876 54970 65900 54972
rect 65956 54970 65962 54972
rect 65716 54918 65718 54970
rect 65898 54918 65900 54970
rect 65654 54916 65660 54918
rect 65716 54916 65740 54918
rect 65796 54916 65820 54918
rect 65876 54916 65900 54918
rect 65956 54916 65962 54918
rect 65654 54896 65962 54916
rect 65654 53884 65962 53904
rect 65654 53882 65660 53884
rect 65716 53882 65740 53884
rect 65796 53882 65820 53884
rect 65876 53882 65900 53884
rect 65956 53882 65962 53884
rect 65716 53830 65718 53882
rect 65898 53830 65900 53882
rect 65654 53828 65660 53830
rect 65716 53828 65740 53830
rect 65796 53828 65820 53830
rect 65876 53828 65900 53830
rect 65956 53828 65962 53830
rect 65654 53808 65962 53828
rect 65654 52796 65962 52816
rect 65654 52794 65660 52796
rect 65716 52794 65740 52796
rect 65796 52794 65820 52796
rect 65876 52794 65900 52796
rect 65956 52794 65962 52796
rect 65716 52742 65718 52794
rect 65898 52742 65900 52794
rect 65654 52740 65660 52742
rect 65716 52740 65740 52742
rect 65796 52740 65820 52742
rect 65876 52740 65900 52742
rect 65956 52740 65962 52742
rect 65654 52720 65962 52740
rect 77404 52018 77432 59366
rect 77392 52012 77444 52018
rect 77392 51954 77444 51960
rect 65654 51708 65962 51728
rect 65654 51706 65660 51708
rect 65716 51706 65740 51708
rect 65796 51706 65820 51708
rect 65876 51706 65900 51708
rect 65956 51706 65962 51708
rect 65716 51654 65718 51706
rect 65898 51654 65900 51706
rect 65654 51652 65660 51654
rect 65716 51652 65740 51654
rect 65796 51652 65820 51654
rect 65876 51652 65900 51654
rect 65956 51652 65962 51654
rect 65654 51632 65962 51652
rect 65654 50620 65962 50640
rect 65654 50618 65660 50620
rect 65716 50618 65740 50620
rect 65796 50618 65820 50620
rect 65876 50618 65900 50620
rect 65956 50618 65962 50620
rect 65716 50566 65718 50618
rect 65898 50566 65900 50618
rect 65654 50564 65660 50566
rect 65716 50564 65740 50566
rect 65796 50564 65820 50566
rect 65876 50564 65900 50566
rect 65956 50564 65962 50566
rect 65654 50544 65962 50564
rect 65654 49532 65962 49552
rect 65654 49530 65660 49532
rect 65716 49530 65740 49532
rect 65796 49530 65820 49532
rect 65876 49530 65900 49532
rect 65956 49530 65962 49532
rect 65716 49478 65718 49530
rect 65898 49478 65900 49530
rect 65654 49476 65660 49478
rect 65716 49476 65740 49478
rect 65796 49476 65820 49478
rect 65876 49476 65900 49478
rect 65956 49476 65962 49478
rect 65654 49456 65962 49476
rect 65654 48444 65962 48464
rect 65654 48442 65660 48444
rect 65716 48442 65740 48444
rect 65796 48442 65820 48444
rect 65876 48442 65900 48444
rect 65956 48442 65962 48444
rect 65716 48390 65718 48442
rect 65898 48390 65900 48442
rect 65654 48388 65660 48390
rect 65716 48388 65740 48390
rect 65796 48388 65820 48390
rect 65876 48388 65900 48390
rect 65956 48388 65962 48390
rect 65654 48368 65962 48388
rect 75828 48272 75880 48278
rect 75828 48214 75880 48220
rect 75840 47705 75868 48214
rect 75826 47696 75882 47705
rect 75826 47631 75882 47640
rect 65654 47356 65962 47376
rect 65654 47354 65660 47356
rect 65716 47354 65740 47356
rect 65796 47354 65820 47356
rect 65876 47354 65900 47356
rect 65956 47354 65962 47356
rect 65716 47302 65718 47354
rect 65898 47302 65900 47354
rect 65654 47300 65660 47302
rect 65716 47300 65740 47302
rect 65796 47300 65820 47302
rect 65876 47300 65900 47302
rect 65956 47300 65962 47302
rect 65654 47280 65962 47300
rect 65654 46268 65962 46288
rect 65654 46266 65660 46268
rect 65716 46266 65740 46268
rect 65796 46266 65820 46268
rect 65876 46266 65900 46268
rect 65956 46266 65962 46268
rect 65716 46214 65718 46266
rect 65898 46214 65900 46266
rect 65654 46212 65660 46214
rect 65716 46212 65740 46214
rect 65796 46212 65820 46214
rect 65876 46212 65900 46214
rect 65956 46212 65962 46214
rect 65654 46192 65962 46212
rect 65654 45180 65962 45200
rect 65654 45178 65660 45180
rect 65716 45178 65740 45180
rect 65796 45178 65820 45180
rect 65876 45178 65900 45180
rect 65956 45178 65962 45180
rect 65716 45126 65718 45178
rect 65898 45126 65900 45178
rect 65654 45124 65660 45126
rect 65716 45124 65740 45126
rect 65796 45124 65820 45126
rect 65876 45124 65900 45126
rect 65956 45124 65962 45126
rect 65654 45104 65962 45124
rect 65654 44092 65962 44112
rect 65654 44090 65660 44092
rect 65716 44090 65740 44092
rect 65796 44090 65820 44092
rect 65876 44090 65900 44092
rect 65956 44090 65962 44092
rect 65716 44038 65718 44090
rect 65898 44038 65900 44090
rect 65654 44036 65660 44038
rect 65716 44036 65740 44038
rect 65796 44036 65820 44038
rect 65876 44036 65900 44038
rect 65956 44036 65962 44038
rect 65654 44016 65962 44036
rect 76564 43784 76616 43790
rect 76564 43726 76616 43732
rect 65654 43004 65962 43024
rect 65654 43002 65660 43004
rect 65716 43002 65740 43004
rect 65796 43002 65820 43004
rect 65876 43002 65900 43004
rect 65956 43002 65962 43004
rect 65716 42950 65718 43002
rect 65898 42950 65900 43002
rect 65654 42948 65660 42950
rect 65716 42948 65740 42950
rect 65796 42948 65820 42950
rect 65876 42948 65900 42950
rect 65956 42948 65962 42950
rect 65654 42928 65962 42948
rect 65654 41916 65962 41936
rect 65654 41914 65660 41916
rect 65716 41914 65740 41916
rect 65796 41914 65820 41916
rect 65876 41914 65900 41916
rect 65956 41914 65962 41916
rect 65716 41862 65718 41914
rect 65898 41862 65900 41914
rect 65654 41860 65660 41862
rect 65716 41860 65740 41862
rect 65796 41860 65820 41862
rect 65876 41860 65900 41862
rect 65956 41860 65962 41862
rect 65654 41840 65962 41860
rect 65654 40828 65962 40848
rect 65654 40826 65660 40828
rect 65716 40826 65740 40828
rect 65796 40826 65820 40828
rect 65876 40826 65900 40828
rect 65956 40826 65962 40828
rect 65716 40774 65718 40826
rect 65898 40774 65900 40826
rect 65654 40772 65660 40774
rect 65716 40772 65740 40774
rect 65796 40772 65820 40774
rect 65876 40772 65900 40774
rect 65956 40772 65962 40774
rect 65654 40752 65962 40772
rect 65654 39740 65962 39760
rect 65654 39738 65660 39740
rect 65716 39738 65740 39740
rect 65796 39738 65820 39740
rect 65876 39738 65900 39740
rect 65956 39738 65962 39740
rect 65716 39686 65718 39738
rect 65898 39686 65900 39738
rect 65654 39684 65660 39686
rect 65716 39684 65740 39686
rect 65796 39684 65820 39686
rect 65876 39684 65900 39686
rect 65956 39684 65962 39686
rect 65654 39664 65962 39684
rect 65654 38652 65962 38672
rect 65654 38650 65660 38652
rect 65716 38650 65740 38652
rect 65796 38650 65820 38652
rect 65876 38650 65900 38652
rect 65956 38650 65962 38652
rect 65716 38598 65718 38650
rect 65898 38598 65900 38650
rect 65654 38596 65660 38598
rect 65716 38596 65740 38598
rect 65796 38596 65820 38598
rect 65876 38596 65900 38598
rect 65956 38596 65962 38598
rect 65654 38576 65962 38596
rect 65654 37564 65962 37584
rect 65654 37562 65660 37564
rect 65716 37562 65740 37564
rect 65796 37562 65820 37564
rect 65876 37562 65900 37564
rect 65956 37562 65962 37564
rect 65716 37510 65718 37562
rect 65898 37510 65900 37562
rect 65654 37508 65660 37510
rect 65716 37508 65740 37510
rect 65796 37508 65820 37510
rect 65876 37508 65900 37510
rect 65956 37508 65962 37510
rect 65654 37488 65962 37508
rect 65654 36476 65962 36496
rect 65654 36474 65660 36476
rect 65716 36474 65740 36476
rect 65796 36474 65820 36476
rect 65876 36474 65900 36476
rect 65956 36474 65962 36476
rect 65716 36422 65718 36474
rect 65898 36422 65900 36474
rect 65654 36420 65660 36422
rect 65716 36420 65740 36422
rect 65796 36420 65820 36422
rect 65876 36420 65900 36422
rect 65956 36420 65962 36422
rect 65654 36400 65962 36420
rect 65654 35388 65962 35408
rect 65654 35386 65660 35388
rect 65716 35386 65740 35388
rect 65796 35386 65820 35388
rect 65876 35386 65900 35388
rect 65956 35386 65962 35388
rect 65716 35334 65718 35386
rect 65898 35334 65900 35386
rect 65654 35332 65660 35334
rect 65716 35332 65740 35334
rect 65796 35332 65820 35334
rect 65876 35332 65900 35334
rect 65956 35332 65962 35334
rect 65654 35312 65962 35332
rect 76576 34678 76604 43726
rect 77576 42628 77628 42634
rect 77576 42570 77628 42576
rect 77484 40520 77536 40526
rect 77484 40462 77536 40468
rect 77496 40186 77524 40462
rect 77484 40180 77536 40186
rect 77484 40122 77536 40128
rect 77588 40118 77616 42570
rect 77576 40112 77628 40118
rect 77576 40054 77628 40060
rect 76564 34672 76616 34678
rect 76564 34614 76616 34620
rect 66628 34604 66680 34610
rect 66628 34546 66680 34552
rect 65654 34300 65962 34320
rect 65654 34298 65660 34300
rect 65716 34298 65740 34300
rect 65796 34298 65820 34300
rect 65876 34298 65900 34300
rect 65956 34298 65962 34300
rect 65716 34246 65718 34298
rect 65898 34246 65900 34298
rect 65654 34244 65660 34246
rect 65716 34244 65740 34246
rect 65796 34244 65820 34246
rect 65876 34244 65900 34246
rect 65956 34244 65962 34246
rect 65654 34224 65962 34244
rect 65654 33212 65962 33232
rect 65654 33210 65660 33212
rect 65716 33210 65740 33212
rect 65796 33210 65820 33212
rect 65876 33210 65900 33212
rect 65956 33210 65962 33212
rect 65716 33158 65718 33210
rect 65898 33158 65900 33210
rect 65654 33156 65660 33158
rect 65716 33156 65740 33158
rect 65796 33156 65820 33158
rect 65876 33156 65900 33158
rect 65956 33156 65962 33158
rect 65654 33136 65962 33156
rect 65654 32124 65962 32144
rect 65654 32122 65660 32124
rect 65716 32122 65740 32124
rect 65796 32122 65820 32124
rect 65876 32122 65900 32124
rect 65956 32122 65962 32124
rect 65716 32070 65718 32122
rect 65898 32070 65900 32122
rect 65654 32068 65660 32070
rect 65716 32068 65740 32070
rect 65796 32068 65820 32070
rect 65876 32068 65900 32070
rect 65956 32068 65962 32070
rect 65654 32048 65962 32068
rect 65654 31036 65962 31056
rect 65654 31034 65660 31036
rect 65716 31034 65740 31036
rect 65796 31034 65820 31036
rect 65876 31034 65900 31036
rect 65956 31034 65962 31036
rect 65716 30982 65718 31034
rect 65898 30982 65900 31034
rect 65654 30980 65660 30982
rect 65716 30980 65740 30982
rect 65796 30980 65820 30982
rect 65876 30980 65900 30982
rect 65956 30980 65962 30982
rect 65654 30960 65962 30980
rect 65654 29948 65962 29968
rect 65654 29946 65660 29948
rect 65716 29946 65740 29948
rect 65796 29946 65820 29948
rect 65876 29946 65900 29948
rect 65956 29946 65962 29948
rect 65716 29894 65718 29946
rect 65898 29894 65900 29946
rect 65654 29892 65660 29894
rect 65716 29892 65740 29894
rect 65796 29892 65820 29894
rect 65876 29892 65900 29894
rect 65956 29892 65962 29894
rect 65654 29872 65962 29892
rect 65654 28860 65962 28880
rect 65654 28858 65660 28860
rect 65716 28858 65740 28860
rect 65796 28858 65820 28860
rect 65876 28858 65900 28860
rect 65956 28858 65962 28860
rect 65716 28806 65718 28858
rect 65898 28806 65900 28858
rect 65654 28804 65660 28806
rect 65716 28804 65740 28806
rect 65796 28804 65820 28806
rect 65876 28804 65900 28806
rect 65956 28804 65962 28806
rect 65654 28784 65962 28804
rect 65654 27772 65962 27792
rect 65654 27770 65660 27772
rect 65716 27770 65740 27772
rect 65796 27770 65820 27772
rect 65876 27770 65900 27772
rect 65956 27770 65962 27772
rect 65716 27718 65718 27770
rect 65898 27718 65900 27770
rect 65654 27716 65660 27718
rect 65716 27716 65740 27718
rect 65796 27716 65820 27718
rect 65876 27716 65900 27718
rect 65956 27716 65962 27718
rect 65654 27696 65962 27716
rect 65654 26684 65962 26704
rect 65654 26682 65660 26684
rect 65716 26682 65740 26684
rect 65796 26682 65820 26684
rect 65876 26682 65900 26684
rect 65956 26682 65962 26684
rect 65716 26630 65718 26682
rect 65898 26630 65900 26682
rect 65654 26628 65660 26630
rect 65716 26628 65740 26630
rect 65796 26628 65820 26630
rect 65876 26628 65900 26630
rect 65956 26628 65962 26630
rect 65654 26608 65962 26628
rect 65654 25596 65962 25616
rect 65654 25594 65660 25596
rect 65716 25594 65740 25596
rect 65796 25594 65820 25596
rect 65876 25594 65900 25596
rect 65956 25594 65962 25596
rect 65716 25542 65718 25594
rect 65898 25542 65900 25594
rect 65654 25540 65660 25542
rect 65716 25540 65740 25542
rect 65796 25540 65820 25542
rect 65876 25540 65900 25542
rect 65956 25540 65962 25542
rect 65654 25520 65962 25540
rect 65654 24508 65962 24528
rect 65654 24506 65660 24508
rect 65716 24506 65740 24508
rect 65796 24506 65820 24508
rect 65876 24506 65900 24508
rect 65956 24506 65962 24508
rect 65716 24454 65718 24506
rect 65898 24454 65900 24506
rect 65654 24452 65660 24454
rect 65716 24452 65740 24454
rect 65796 24452 65820 24454
rect 65876 24452 65900 24454
rect 65956 24452 65962 24454
rect 65654 24432 65962 24452
rect 65654 23420 65962 23440
rect 65654 23418 65660 23420
rect 65716 23418 65740 23420
rect 65796 23418 65820 23420
rect 65876 23418 65900 23420
rect 65956 23418 65962 23420
rect 65716 23366 65718 23418
rect 65898 23366 65900 23418
rect 65654 23364 65660 23366
rect 65716 23364 65740 23366
rect 65796 23364 65820 23366
rect 65876 23364 65900 23366
rect 65956 23364 65962 23366
rect 65654 23344 65962 23364
rect 65654 22332 65962 22352
rect 65654 22330 65660 22332
rect 65716 22330 65740 22332
rect 65796 22330 65820 22332
rect 65876 22330 65900 22332
rect 65956 22330 65962 22332
rect 65716 22278 65718 22330
rect 65898 22278 65900 22330
rect 65654 22276 65660 22278
rect 65716 22276 65740 22278
rect 65796 22276 65820 22278
rect 65876 22276 65900 22278
rect 65956 22276 65962 22278
rect 65654 22256 65962 22276
rect 65654 21244 65962 21264
rect 65654 21242 65660 21244
rect 65716 21242 65740 21244
rect 65796 21242 65820 21244
rect 65876 21242 65900 21244
rect 65956 21242 65962 21244
rect 65716 21190 65718 21242
rect 65898 21190 65900 21242
rect 65654 21188 65660 21190
rect 65716 21188 65740 21190
rect 65796 21188 65820 21190
rect 65876 21188 65900 21190
rect 65956 21188 65962 21190
rect 65654 21168 65962 21188
rect 65654 20156 65962 20176
rect 65654 20154 65660 20156
rect 65716 20154 65740 20156
rect 65796 20154 65820 20156
rect 65876 20154 65900 20156
rect 65956 20154 65962 20156
rect 65716 20102 65718 20154
rect 65898 20102 65900 20154
rect 65654 20100 65660 20102
rect 65716 20100 65740 20102
rect 65796 20100 65820 20102
rect 65876 20100 65900 20102
rect 65956 20100 65962 20102
rect 65654 20080 65962 20100
rect 65654 19068 65962 19088
rect 65654 19066 65660 19068
rect 65716 19066 65740 19068
rect 65796 19066 65820 19068
rect 65876 19066 65900 19068
rect 65956 19066 65962 19068
rect 65716 19014 65718 19066
rect 65898 19014 65900 19066
rect 65654 19012 65660 19014
rect 65716 19012 65740 19014
rect 65796 19012 65820 19014
rect 65876 19012 65900 19014
rect 65956 19012 65962 19014
rect 65654 18992 65962 19012
rect 65654 17980 65962 18000
rect 65654 17978 65660 17980
rect 65716 17978 65740 17980
rect 65796 17978 65820 17980
rect 65876 17978 65900 17980
rect 65956 17978 65962 17980
rect 65716 17926 65718 17978
rect 65898 17926 65900 17978
rect 65654 17924 65660 17926
rect 65716 17924 65740 17926
rect 65796 17924 65820 17926
rect 65876 17924 65900 17926
rect 65956 17924 65962 17926
rect 65654 17904 65962 17924
rect 65654 16892 65962 16912
rect 65654 16890 65660 16892
rect 65716 16890 65740 16892
rect 65796 16890 65820 16892
rect 65876 16890 65900 16892
rect 65956 16890 65962 16892
rect 65716 16838 65718 16890
rect 65898 16838 65900 16890
rect 65654 16836 65660 16838
rect 65716 16836 65740 16838
rect 65796 16836 65820 16838
rect 65876 16836 65900 16838
rect 65956 16836 65962 16838
rect 65654 16816 65962 16836
rect 63040 16584 63092 16590
rect 41156 16546 41276 16574
rect 41144 3392 41196 3398
rect 41144 3334 41196 3340
rect 41052 2576 41104 2582
rect 40880 2502 41000 2530
rect 41052 2518 41104 2524
rect 41156 2514 41184 3334
rect 41248 2990 41276 16546
rect 63040 16526 63092 16532
rect 50294 16348 50602 16368
rect 50294 16346 50300 16348
rect 50356 16346 50380 16348
rect 50436 16346 50460 16348
rect 50516 16346 50540 16348
rect 50596 16346 50602 16348
rect 50356 16294 50358 16346
rect 50538 16294 50540 16346
rect 50294 16292 50300 16294
rect 50356 16292 50380 16294
rect 50436 16292 50460 16294
rect 50516 16292 50540 16294
rect 50596 16292 50602 16294
rect 50294 16272 50602 16292
rect 65654 15804 65962 15824
rect 65654 15802 65660 15804
rect 65716 15802 65740 15804
rect 65796 15802 65820 15804
rect 65876 15802 65900 15804
rect 65956 15802 65962 15804
rect 65716 15750 65718 15802
rect 65898 15750 65900 15802
rect 65654 15748 65660 15750
rect 65716 15748 65740 15750
rect 65796 15748 65820 15750
rect 65876 15748 65900 15750
rect 65956 15748 65962 15750
rect 65654 15728 65962 15748
rect 50294 15260 50602 15280
rect 50294 15258 50300 15260
rect 50356 15258 50380 15260
rect 50436 15258 50460 15260
rect 50516 15258 50540 15260
rect 50596 15258 50602 15260
rect 50356 15206 50358 15258
rect 50538 15206 50540 15258
rect 50294 15204 50300 15206
rect 50356 15204 50380 15206
rect 50436 15204 50460 15206
rect 50516 15204 50540 15206
rect 50596 15204 50602 15206
rect 50294 15184 50602 15204
rect 65654 14716 65962 14736
rect 65654 14714 65660 14716
rect 65716 14714 65740 14716
rect 65796 14714 65820 14716
rect 65876 14714 65900 14716
rect 65956 14714 65962 14716
rect 65716 14662 65718 14714
rect 65898 14662 65900 14714
rect 65654 14660 65660 14662
rect 65716 14660 65740 14662
rect 65796 14660 65820 14662
rect 65876 14660 65900 14662
rect 65956 14660 65962 14662
rect 65654 14640 65962 14660
rect 50294 14172 50602 14192
rect 50294 14170 50300 14172
rect 50356 14170 50380 14172
rect 50436 14170 50460 14172
rect 50516 14170 50540 14172
rect 50596 14170 50602 14172
rect 50356 14118 50358 14170
rect 50538 14118 50540 14170
rect 50294 14116 50300 14118
rect 50356 14116 50380 14118
rect 50436 14116 50460 14118
rect 50516 14116 50540 14118
rect 50596 14116 50602 14118
rect 50294 14096 50602 14116
rect 65654 13628 65962 13648
rect 65654 13626 65660 13628
rect 65716 13626 65740 13628
rect 65796 13626 65820 13628
rect 65876 13626 65900 13628
rect 65956 13626 65962 13628
rect 65716 13574 65718 13626
rect 65898 13574 65900 13626
rect 65654 13572 65660 13574
rect 65716 13572 65740 13574
rect 65796 13572 65820 13574
rect 65876 13572 65900 13574
rect 65956 13572 65962 13574
rect 65654 13552 65962 13572
rect 50294 13084 50602 13104
rect 50294 13082 50300 13084
rect 50356 13082 50380 13084
rect 50436 13082 50460 13084
rect 50516 13082 50540 13084
rect 50596 13082 50602 13084
rect 50356 13030 50358 13082
rect 50538 13030 50540 13082
rect 50294 13028 50300 13030
rect 50356 13028 50380 13030
rect 50436 13028 50460 13030
rect 50516 13028 50540 13030
rect 50596 13028 50602 13030
rect 50294 13008 50602 13028
rect 65654 12540 65962 12560
rect 65654 12538 65660 12540
rect 65716 12538 65740 12540
rect 65796 12538 65820 12540
rect 65876 12538 65900 12540
rect 65956 12538 65962 12540
rect 65716 12486 65718 12538
rect 65898 12486 65900 12538
rect 65654 12484 65660 12486
rect 65716 12484 65740 12486
rect 65796 12484 65820 12486
rect 65876 12484 65900 12486
rect 65956 12484 65962 12486
rect 65654 12464 65962 12484
rect 50294 11996 50602 12016
rect 50294 11994 50300 11996
rect 50356 11994 50380 11996
rect 50436 11994 50460 11996
rect 50516 11994 50540 11996
rect 50596 11994 50602 11996
rect 50356 11942 50358 11994
rect 50538 11942 50540 11994
rect 50294 11940 50300 11942
rect 50356 11940 50380 11942
rect 50436 11940 50460 11942
rect 50516 11940 50540 11942
rect 50596 11940 50602 11942
rect 50294 11920 50602 11940
rect 65654 11452 65962 11472
rect 65654 11450 65660 11452
rect 65716 11450 65740 11452
rect 65796 11450 65820 11452
rect 65876 11450 65900 11452
rect 65956 11450 65962 11452
rect 65716 11398 65718 11450
rect 65898 11398 65900 11450
rect 65654 11396 65660 11398
rect 65716 11396 65740 11398
rect 65796 11396 65820 11398
rect 65876 11396 65900 11398
rect 65956 11396 65962 11398
rect 65654 11376 65962 11396
rect 50294 10908 50602 10928
rect 50294 10906 50300 10908
rect 50356 10906 50380 10908
rect 50436 10906 50460 10908
rect 50516 10906 50540 10908
rect 50596 10906 50602 10908
rect 50356 10854 50358 10906
rect 50538 10854 50540 10906
rect 50294 10852 50300 10854
rect 50356 10852 50380 10854
rect 50436 10852 50460 10854
rect 50516 10852 50540 10854
rect 50596 10852 50602 10854
rect 50294 10832 50602 10852
rect 65654 10364 65962 10384
rect 65654 10362 65660 10364
rect 65716 10362 65740 10364
rect 65796 10362 65820 10364
rect 65876 10362 65900 10364
rect 65956 10362 65962 10364
rect 65716 10310 65718 10362
rect 65898 10310 65900 10362
rect 65654 10308 65660 10310
rect 65716 10308 65740 10310
rect 65796 10308 65820 10310
rect 65876 10308 65900 10310
rect 65956 10308 65962 10310
rect 65654 10288 65962 10308
rect 50294 9820 50602 9840
rect 50294 9818 50300 9820
rect 50356 9818 50380 9820
rect 50436 9818 50460 9820
rect 50516 9818 50540 9820
rect 50596 9818 50602 9820
rect 50356 9766 50358 9818
rect 50538 9766 50540 9818
rect 50294 9764 50300 9766
rect 50356 9764 50380 9766
rect 50436 9764 50460 9766
rect 50516 9764 50540 9766
rect 50596 9764 50602 9766
rect 50294 9744 50602 9764
rect 65654 9276 65962 9296
rect 65654 9274 65660 9276
rect 65716 9274 65740 9276
rect 65796 9274 65820 9276
rect 65876 9274 65900 9276
rect 65956 9274 65962 9276
rect 65716 9222 65718 9274
rect 65898 9222 65900 9274
rect 65654 9220 65660 9222
rect 65716 9220 65740 9222
rect 65796 9220 65820 9222
rect 65876 9220 65900 9222
rect 65956 9220 65962 9222
rect 65654 9200 65962 9220
rect 50294 8732 50602 8752
rect 50294 8730 50300 8732
rect 50356 8730 50380 8732
rect 50436 8730 50460 8732
rect 50516 8730 50540 8732
rect 50596 8730 50602 8732
rect 50356 8678 50358 8730
rect 50538 8678 50540 8730
rect 50294 8676 50300 8678
rect 50356 8676 50380 8678
rect 50436 8676 50460 8678
rect 50516 8676 50540 8678
rect 50596 8676 50602 8678
rect 50294 8656 50602 8676
rect 65654 8188 65962 8208
rect 65654 8186 65660 8188
rect 65716 8186 65740 8188
rect 65796 8186 65820 8188
rect 65876 8186 65900 8188
rect 65956 8186 65962 8188
rect 65716 8134 65718 8186
rect 65898 8134 65900 8186
rect 65654 8132 65660 8134
rect 65716 8132 65740 8134
rect 65796 8132 65820 8134
rect 65876 8132 65900 8134
rect 65956 8132 65962 8134
rect 65654 8112 65962 8132
rect 50294 7644 50602 7664
rect 50294 7642 50300 7644
rect 50356 7642 50380 7644
rect 50436 7642 50460 7644
rect 50516 7642 50540 7644
rect 50596 7642 50602 7644
rect 50356 7590 50358 7642
rect 50538 7590 50540 7642
rect 50294 7588 50300 7590
rect 50356 7588 50380 7590
rect 50436 7588 50460 7590
rect 50516 7588 50540 7590
rect 50596 7588 50602 7590
rect 50294 7568 50602 7588
rect 65654 7100 65962 7120
rect 65654 7098 65660 7100
rect 65716 7098 65740 7100
rect 65796 7098 65820 7100
rect 65876 7098 65900 7100
rect 65956 7098 65962 7100
rect 65716 7046 65718 7098
rect 65898 7046 65900 7098
rect 65654 7044 65660 7046
rect 65716 7044 65740 7046
rect 65796 7044 65820 7046
rect 65876 7044 65900 7046
rect 65956 7044 65962 7046
rect 65654 7024 65962 7044
rect 50294 6556 50602 6576
rect 50294 6554 50300 6556
rect 50356 6554 50380 6556
rect 50436 6554 50460 6556
rect 50516 6554 50540 6556
rect 50596 6554 50602 6556
rect 50356 6502 50358 6554
rect 50538 6502 50540 6554
rect 50294 6500 50300 6502
rect 50356 6500 50380 6502
rect 50436 6500 50460 6502
rect 50516 6500 50540 6502
rect 50596 6500 50602 6502
rect 50294 6480 50602 6500
rect 65654 6012 65962 6032
rect 65654 6010 65660 6012
rect 65716 6010 65740 6012
rect 65796 6010 65820 6012
rect 65876 6010 65900 6012
rect 65956 6010 65962 6012
rect 65716 5958 65718 6010
rect 65898 5958 65900 6010
rect 65654 5956 65660 5958
rect 65716 5956 65740 5958
rect 65796 5956 65820 5958
rect 65876 5956 65900 5958
rect 65956 5956 65962 5958
rect 65654 5936 65962 5956
rect 50294 5468 50602 5488
rect 50294 5466 50300 5468
rect 50356 5466 50380 5468
rect 50436 5466 50460 5468
rect 50516 5466 50540 5468
rect 50596 5466 50602 5468
rect 50356 5414 50358 5466
rect 50538 5414 50540 5466
rect 50294 5412 50300 5414
rect 50356 5412 50380 5414
rect 50436 5412 50460 5414
rect 50516 5412 50540 5414
rect 50596 5412 50602 5414
rect 50294 5392 50602 5412
rect 65654 4924 65962 4944
rect 65654 4922 65660 4924
rect 65716 4922 65740 4924
rect 65796 4922 65820 4924
rect 65876 4922 65900 4924
rect 65956 4922 65962 4924
rect 65716 4870 65718 4922
rect 65898 4870 65900 4922
rect 65654 4868 65660 4870
rect 65716 4868 65740 4870
rect 65796 4868 65820 4870
rect 65876 4868 65900 4870
rect 65956 4868 65962 4870
rect 65654 4848 65962 4868
rect 50294 4380 50602 4400
rect 50294 4378 50300 4380
rect 50356 4378 50380 4380
rect 50436 4378 50460 4380
rect 50516 4378 50540 4380
rect 50596 4378 50602 4380
rect 50356 4326 50358 4378
rect 50538 4326 50540 4378
rect 50294 4324 50300 4326
rect 50356 4324 50380 4326
rect 50436 4324 50460 4326
rect 50516 4324 50540 4326
rect 50596 4324 50602 4326
rect 50294 4304 50602 4324
rect 65654 3836 65962 3856
rect 65654 3834 65660 3836
rect 65716 3834 65740 3836
rect 65796 3834 65820 3836
rect 65876 3834 65900 3836
rect 65956 3834 65962 3836
rect 65716 3782 65718 3834
rect 65898 3782 65900 3834
rect 65654 3780 65660 3782
rect 65716 3780 65740 3782
rect 65796 3780 65820 3782
rect 65876 3780 65900 3782
rect 65956 3780 65962 3782
rect 65654 3760 65962 3780
rect 43904 3528 43956 3534
rect 43904 3470 43956 3476
rect 41696 3392 41748 3398
rect 41696 3334 41748 3340
rect 41236 2984 41288 2990
rect 41236 2926 41288 2932
rect 40972 2310 41000 2502
rect 41144 2508 41196 2514
rect 41144 2450 41196 2456
rect 41708 2446 41736 3334
rect 43916 2650 43944 3470
rect 57980 3460 58032 3466
rect 57980 3402 58032 3408
rect 50294 3292 50602 3312
rect 50294 3290 50300 3292
rect 50356 3290 50380 3292
rect 50436 3290 50460 3292
rect 50516 3290 50540 3292
rect 50596 3290 50602 3292
rect 50356 3238 50358 3290
rect 50538 3238 50540 3290
rect 50294 3236 50300 3238
rect 50356 3236 50380 3238
rect 50436 3236 50460 3238
rect 50516 3236 50540 3238
rect 50596 3236 50602 3238
rect 50294 3216 50602 3236
rect 43904 2644 43956 2650
rect 43904 2586 43956 2592
rect 55772 2644 55824 2650
rect 55772 2586 55824 2592
rect 50620 2576 50672 2582
rect 50620 2518 50672 2524
rect 41696 2440 41748 2446
rect 41696 2382 41748 2388
rect 44456 2440 44508 2446
rect 44456 2382 44508 2388
rect 47676 2440 47728 2446
rect 47676 2382 47728 2388
rect 40592 2304 40644 2310
rect 40592 2246 40644 2252
rect 40960 2304 41012 2310
rect 40960 2246 41012 2252
rect 39948 1964 40000 1970
rect 39948 1906 40000 1912
rect 40604 800 40632 2246
rect 44468 800 44496 2382
rect 47688 800 47716 2382
rect 50632 2310 50660 2518
rect 55784 2446 55812 2586
rect 51540 2440 51592 2446
rect 51540 2382 51592 2388
rect 55404 2440 55456 2446
rect 55404 2382 55456 2388
rect 55772 2440 55824 2446
rect 55772 2382 55824 2388
rect 50620 2304 50672 2310
rect 50620 2246 50672 2252
rect 50294 2204 50602 2224
rect 50294 2202 50300 2204
rect 50356 2202 50380 2204
rect 50436 2202 50460 2204
rect 50516 2202 50540 2204
rect 50596 2202 50602 2204
rect 50356 2150 50358 2202
rect 50538 2150 50540 2202
rect 50294 2148 50300 2150
rect 50356 2148 50380 2150
rect 50436 2148 50460 2150
rect 50516 2148 50540 2150
rect 50596 2148 50602 2150
rect 50294 2128 50602 2148
rect 51552 800 51580 2382
rect 51908 2372 51960 2378
rect 51908 2314 51960 2320
rect 51920 1970 51948 2314
rect 51908 1964 51960 1970
rect 51908 1906 51960 1912
rect 55416 800 55444 2382
rect 57992 2378 58020 3402
rect 65654 2748 65962 2768
rect 65654 2746 65660 2748
rect 65716 2746 65740 2748
rect 65796 2746 65820 2748
rect 65876 2746 65900 2748
rect 65956 2746 65962 2748
rect 65716 2694 65718 2746
rect 65898 2694 65900 2746
rect 65654 2692 65660 2694
rect 65716 2692 65740 2694
rect 65796 2692 65820 2694
rect 65876 2692 65900 2694
rect 65956 2692 65962 2694
rect 65654 2672 65962 2692
rect 66640 2650 66668 34546
rect 77208 12844 77260 12850
rect 77208 12786 77260 12792
rect 77220 12345 77248 12786
rect 77206 12336 77262 12345
rect 77206 12271 77262 12280
rect 66628 2644 66680 2650
rect 66628 2586 66680 2592
rect 59268 2440 59320 2446
rect 59268 2382 59320 2388
rect 62488 2440 62540 2446
rect 62488 2382 62540 2388
rect 66352 2440 66404 2446
rect 66352 2382 66404 2388
rect 70216 2440 70268 2446
rect 70216 2382 70268 2388
rect 77300 2440 77352 2446
rect 77300 2382 77352 2388
rect 57980 2372 58032 2378
rect 57980 2314 58032 2320
rect 59280 800 59308 2382
rect 62500 800 62528 2382
rect 63868 2372 63920 2378
rect 63868 2314 63920 2320
rect 63880 2038 63908 2314
rect 63868 2032 63920 2038
rect 63868 1974 63920 1980
rect 66364 800 66392 2382
rect 70228 800 70256 2382
rect 74080 2304 74132 2310
rect 74080 2246 74132 2252
rect 74092 800 74120 2246
rect 77312 800 77340 2382
rect 77588 1902 77616 40054
rect 77680 12918 77708 70926
rect 77772 60314 77800 110706
rect 77852 110560 77904 110566
rect 77852 110502 77904 110508
rect 77864 110265 77892 110502
rect 77850 110256 77906 110265
rect 77850 110191 77906 110200
rect 77852 106208 77904 106214
rect 77850 106176 77852 106185
rect 77904 106176 77906 106185
rect 77850 106111 77906 106120
rect 77944 103760 77996 103766
rect 77944 103702 77996 103708
rect 77852 102944 77904 102950
rect 77852 102886 77904 102892
rect 77864 102785 77892 102886
rect 77850 102776 77906 102785
rect 77850 102711 77906 102720
rect 77850 98696 77906 98705
rect 77850 98631 77852 98640
rect 77904 98631 77906 98640
rect 77852 98602 77904 98608
rect 77956 94926 77984 103702
rect 78048 103630 78076 113146
rect 78036 103624 78088 103630
rect 78036 103566 78088 103572
rect 78128 98796 78180 98802
rect 78128 98738 78180 98744
rect 77944 94920 77996 94926
rect 77944 94862 77996 94868
rect 78036 94784 78088 94790
rect 78036 94726 78088 94732
rect 78048 94625 78076 94726
rect 78034 94616 78090 94625
rect 78034 94551 78090 94560
rect 77942 90536 77998 90545
rect 77942 90471 77944 90480
rect 77996 90471 77998 90480
rect 77944 90442 77996 90448
rect 77944 87236 77996 87242
rect 77944 87178 77996 87184
rect 77956 87145 77984 87178
rect 77942 87136 77998 87145
rect 77942 87071 77998 87080
rect 77852 83360 77904 83366
rect 77852 83302 77904 83308
rect 77864 83065 77892 83302
rect 77850 83056 77906 83065
rect 77850 82991 77906 83000
rect 77944 75336 77996 75342
rect 77944 75278 77996 75284
rect 77850 71496 77906 71505
rect 77850 71431 77852 71440
rect 77904 71431 77906 71440
rect 77852 71402 77904 71408
rect 77956 69766 77984 75278
rect 78036 75200 78088 75206
rect 78036 75142 78088 75148
rect 78048 74905 78076 75142
rect 78034 74896 78090 74905
rect 78034 74831 78090 74840
rect 77944 69760 77996 69766
rect 77944 69702 77996 69708
rect 77944 67652 77996 67658
rect 77944 67594 77996 67600
rect 77852 67584 77904 67590
rect 77852 67526 77904 67532
rect 77864 64870 77892 67526
rect 77956 67425 77984 67594
rect 77942 67416 77998 67425
rect 77942 67351 77998 67360
rect 77852 64864 77904 64870
rect 77852 64806 77904 64812
rect 78034 63336 78090 63345
rect 78034 63271 78090 63280
rect 78048 63238 78076 63271
rect 78036 63232 78088 63238
rect 78036 63174 78088 63180
rect 77760 60308 77812 60314
rect 77760 60250 77812 60256
rect 77760 60036 77812 60042
rect 77760 59978 77812 59984
rect 77772 59770 77800 59978
rect 77760 59764 77812 59770
rect 77760 59706 77812 59712
rect 77944 59628 77996 59634
rect 77944 59570 77996 59576
rect 77956 59265 77984 59570
rect 77942 59256 77998 59265
rect 77942 59191 77998 59200
rect 77760 56364 77812 56370
rect 77760 56306 77812 56312
rect 77772 42770 77800 56306
rect 77852 56160 77904 56166
rect 77852 56102 77904 56108
rect 77864 55865 77892 56102
rect 77850 55856 77906 55865
rect 77850 55791 77906 55800
rect 77852 51808 77904 51814
rect 77850 51776 77852 51785
rect 77904 51776 77906 51785
rect 77850 51711 77906 51720
rect 78036 43648 78088 43654
rect 78034 43616 78036 43625
rect 78088 43616 78090 43625
rect 78034 43551 78090 43560
rect 77760 42764 77812 42770
rect 77760 42706 77812 42712
rect 78036 40384 78088 40390
rect 78036 40326 78088 40332
rect 78048 40225 78076 40326
rect 78034 40216 78090 40225
rect 78034 40151 78090 40160
rect 77852 36168 77904 36174
rect 77852 36110 77904 36116
rect 78034 36136 78090 36145
rect 77864 33114 77892 36110
rect 78034 36071 78090 36080
rect 78048 36038 78076 36071
rect 78036 36032 78088 36038
rect 78036 35974 78088 35980
rect 77852 33108 77904 33114
rect 77852 33050 77904 33056
rect 78036 32904 78088 32910
rect 78036 32846 78088 32852
rect 77760 32428 77812 32434
rect 77760 32370 77812 32376
rect 77772 32065 77800 32370
rect 77852 32224 77904 32230
rect 77852 32166 77904 32172
rect 77758 32056 77814 32065
rect 77758 31991 77814 32000
rect 77864 25906 77892 32166
rect 78048 28218 78076 32846
rect 78036 28212 78088 28218
rect 78036 28154 78088 28160
rect 77944 28076 77996 28082
rect 77944 28018 77996 28024
rect 77956 27985 77984 28018
rect 77942 27976 77998 27985
rect 77942 27911 77998 27920
rect 77852 25900 77904 25906
rect 77852 25842 77904 25848
rect 77852 24608 77904 24614
rect 77850 24576 77852 24585
rect 77904 24576 77906 24585
rect 77850 24511 77906 24520
rect 77760 20936 77812 20942
rect 77760 20878 77812 20884
rect 77668 12912 77720 12918
rect 77668 12854 77720 12860
rect 77772 12102 77800 20878
rect 78036 20800 78088 20806
rect 78036 20742 78088 20748
rect 78048 20505 78076 20742
rect 78034 20496 78090 20505
rect 78034 20431 78090 20440
rect 78036 16448 78088 16454
rect 78034 16416 78036 16425
rect 78088 16416 78090 16425
rect 78034 16351 78090 16360
rect 77760 12096 77812 12102
rect 77760 12038 77812 12044
rect 78140 10130 78168 98738
rect 78128 10124 78180 10130
rect 78128 10066 78180 10072
rect 77944 10056 77996 10062
rect 77944 9998 77996 10004
rect 77956 6914 77984 9998
rect 78034 8936 78090 8945
rect 78034 8871 78090 8880
rect 78048 8838 78076 8871
rect 78036 8832 78088 8838
rect 78036 8774 78088 8780
rect 77956 6886 78076 6914
rect 77668 5228 77720 5234
rect 77668 5170 77720 5176
rect 77680 4826 77708 5170
rect 77852 5024 77904 5030
rect 77852 4966 77904 4972
rect 77864 4865 77892 4966
rect 77850 4856 77906 4865
rect 77668 4820 77720 4826
rect 77850 4791 77906 4800
rect 77668 4762 77720 4768
rect 78048 4622 78076 6886
rect 78036 4616 78088 4622
rect 78036 4558 78088 4564
rect 77668 3052 77720 3058
rect 77668 2994 77720 3000
rect 77576 1896 77628 1902
rect 77576 1838 77628 1844
rect 18 0 74 800
rect 3238 0 3294 800
rect 7102 0 7158 800
rect 10966 0 11022 800
rect 14830 0 14886 800
rect 18050 0 18106 800
rect 21914 0 21970 800
rect 25778 0 25834 800
rect 29642 0 29698 800
rect 32862 0 32918 800
rect 36726 0 36782 800
rect 40590 0 40646 800
rect 44454 0 44510 800
rect 47674 0 47730 800
rect 51538 0 51594 800
rect 55402 0 55458 800
rect 59266 0 59322 800
rect 62486 0 62542 800
rect 66350 0 66406 800
rect 70214 0 70270 800
rect 74078 0 74134 800
rect 77298 0 77354 800
rect 77680 785 77708 2994
rect 78048 2514 78076 4558
rect 78036 2508 78088 2514
rect 78036 2450 78088 2456
rect 77666 776 77722 785
rect 77666 711 77722 720
<< via2 >>
rect 1858 117000 1914 117056
rect 1398 105440 1454 105496
rect 1398 101396 1400 101416
rect 1400 101396 1452 101416
rect 1452 101396 1454 101416
rect 1398 101360 1454 101396
rect 1398 97280 1454 97336
rect 1582 112920 1638 112976
rect 1858 109520 1914 109576
rect 1582 93880 1638 93936
rect 1490 89800 1546 89856
rect 1582 85720 1638 85776
rect 1398 81640 1454 81696
rect 1582 78240 1638 78296
rect 1582 74160 1638 74216
rect 1582 70080 1638 70136
rect 1582 66020 1638 66056
rect 1582 66000 1584 66020
rect 1584 66000 1636 66020
rect 1636 66000 1638 66020
rect 1582 62636 1584 62656
rect 1584 62636 1636 62656
rect 1636 62636 1638 62656
rect 1582 62600 1638 62636
rect 1582 58520 1638 58576
rect 4220 116986 4276 116988
rect 4300 116986 4356 116988
rect 4380 116986 4436 116988
rect 4460 116986 4516 116988
rect 4220 116934 4266 116986
rect 4266 116934 4276 116986
rect 4300 116934 4330 116986
rect 4330 116934 4342 116986
rect 4342 116934 4356 116986
rect 4380 116934 4394 116986
rect 4394 116934 4406 116986
rect 4406 116934 4436 116986
rect 4460 116934 4470 116986
rect 4470 116934 4516 116986
rect 4220 116932 4276 116934
rect 4300 116932 4356 116934
rect 4380 116932 4436 116934
rect 4460 116932 4516 116934
rect 4220 115898 4276 115900
rect 4300 115898 4356 115900
rect 4380 115898 4436 115900
rect 4460 115898 4516 115900
rect 4220 115846 4266 115898
rect 4266 115846 4276 115898
rect 4300 115846 4330 115898
rect 4330 115846 4342 115898
rect 4342 115846 4356 115898
rect 4380 115846 4394 115898
rect 4394 115846 4406 115898
rect 4406 115846 4436 115898
rect 4460 115846 4470 115898
rect 4470 115846 4516 115898
rect 4220 115844 4276 115846
rect 4300 115844 4356 115846
rect 4380 115844 4436 115846
rect 4460 115844 4516 115846
rect 4220 114810 4276 114812
rect 4300 114810 4356 114812
rect 4380 114810 4436 114812
rect 4460 114810 4516 114812
rect 4220 114758 4266 114810
rect 4266 114758 4276 114810
rect 4300 114758 4330 114810
rect 4330 114758 4342 114810
rect 4342 114758 4356 114810
rect 4380 114758 4394 114810
rect 4394 114758 4406 114810
rect 4406 114758 4436 114810
rect 4460 114758 4470 114810
rect 4470 114758 4516 114810
rect 4220 114756 4276 114758
rect 4300 114756 4356 114758
rect 4380 114756 4436 114758
rect 4460 114756 4516 114758
rect 4220 113722 4276 113724
rect 4300 113722 4356 113724
rect 4380 113722 4436 113724
rect 4460 113722 4516 113724
rect 4220 113670 4266 113722
rect 4266 113670 4276 113722
rect 4300 113670 4330 113722
rect 4330 113670 4342 113722
rect 4342 113670 4356 113722
rect 4380 113670 4394 113722
rect 4394 113670 4406 113722
rect 4406 113670 4436 113722
rect 4460 113670 4470 113722
rect 4470 113670 4516 113722
rect 4220 113668 4276 113670
rect 4300 113668 4356 113670
rect 4380 113668 4436 113670
rect 4460 113668 4516 113670
rect 4220 112634 4276 112636
rect 4300 112634 4356 112636
rect 4380 112634 4436 112636
rect 4460 112634 4516 112636
rect 4220 112582 4266 112634
rect 4266 112582 4276 112634
rect 4300 112582 4330 112634
rect 4330 112582 4342 112634
rect 4342 112582 4356 112634
rect 4380 112582 4394 112634
rect 4394 112582 4406 112634
rect 4406 112582 4436 112634
rect 4460 112582 4470 112634
rect 4470 112582 4516 112634
rect 4220 112580 4276 112582
rect 4300 112580 4356 112582
rect 4380 112580 4436 112582
rect 4460 112580 4516 112582
rect 4220 111546 4276 111548
rect 4300 111546 4356 111548
rect 4380 111546 4436 111548
rect 4460 111546 4516 111548
rect 4220 111494 4266 111546
rect 4266 111494 4276 111546
rect 4300 111494 4330 111546
rect 4330 111494 4342 111546
rect 4342 111494 4356 111546
rect 4380 111494 4394 111546
rect 4394 111494 4406 111546
rect 4406 111494 4436 111546
rect 4460 111494 4470 111546
rect 4470 111494 4516 111546
rect 4220 111492 4276 111494
rect 4300 111492 4356 111494
rect 4380 111492 4436 111494
rect 4460 111492 4516 111494
rect 4220 110458 4276 110460
rect 4300 110458 4356 110460
rect 4380 110458 4436 110460
rect 4460 110458 4516 110460
rect 4220 110406 4266 110458
rect 4266 110406 4276 110458
rect 4300 110406 4330 110458
rect 4330 110406 4342 110458
rect 4342 110406 4356 110458
rect 4380 110406 4394 110458
rect 4394 110406 4406 110458
rect 4406 110406 4436 110458
rect 4460 110406 4470 110458
rect 4470 110406 4516 110458
rect 4220 110404 4276 110406
rect 4300 110404 4356 110406
rect 4380 110404 4436 110406
rect 4460 110404 4516 110406
rect 4220 109370 4276 109372
rect 4300 109370 4356 109372
rect 4380 109370 4436 109372
rect 4460 109370 4516 109372
rect 4220 109318 4266 109370
rect 4266 109318 4276 109370
rect 4300 109318 4330 109370
rect 4330 109318 4342 109370
rect 4342 109318 4356 109370
rect 4380 109318 4394 109370
rect 4394 109318 4406 109370
rect 4406 109318 4436 109370
rect 4460 109318 4470 109370
rect 4470 109318 4516 109370
rect 4220 109316 4276 109318
rect 4300 109316 4356 109318
rect 4380 109316 4436 109318
rect 4460 109316 4516 109318
rect 4220 108282 4276 108284
rect 4300 108282 4356 108284
rect 4380 108282 4436 108284
rect 4460 108282 4516 108284
rect 4220 108230 4266 108282
rect 4266 108230 4276 108282
rect 4300 108230 4330 108282
rect 4330 108230 4342 108282
rect 4342 108230 4356 108282
rect 4380 108230 4394 108282
rect 4394 108230 4406 108282
rect 4406 108230 4436 108282
rect 4460 108230 4470 108282
rect 4470 108230 4516 108282
rect 4220 108228 4276 108230
rect 4300 108228 4356 108230
rect 4380 108228 4436 108230
rect 4460 108228 4516 108230
rect 4220 107194 4276 107196
rect 4300 107194 4356 107196
rect 4380 107194 4436 107196
rect 4460 107194 4516 107196
rect 4220 107142 4266 107194
rect 4266 107142 4276 107194
rect 4300 107142 4330 107194
rect 4330 107142 4342 107194
rect 4342 107142 4356 107194
rect 4380 107142 4394 107194
rect 4394 107142 4406 107194
rect 4406 107142 4436 107194
rect 4460 107142 4470 107194
rect 4470 107142 4516 107194
rect 4220 107140 4276 107142
rect 4300 107140 4356 107142
rect 4380 107140 4436 107142
rect 4460 107140 4516 107142
rect 4220 106106 4276 106108
rect 4300 106106 4356 106108
rect 4380 106106 4436 106108
rect 4460 106106 4516 106108
rect 4220 106054 4266 106106
rect 4266 106054 4276 106106
rect 4300 106054 4330 106106
rect 4330 106054 4342 106106
rect 4342 106054 4356 106106
rect 4380 106054 4394 106106
rect 4394 106054 4406 106106
rect 4406 106054 4436 106106
rect 4460 106054 4470 106106
rect 4470 106054 4516 106106
rect 4220 106052 4276 106054
rect 4300 106052 4356 106054
rect 4380 106052 4436 106054
rect 4460 106052 4516 106054
rect 4220 105018 4276 105020
rect 4300 105018 4356 105020
rect 4380 105018 4436 105020
rect 4460 105018 4516 105020
rect 4220 104966 4266 105018
rect 4266 104966 4276 105018
rect 4300 104966 4330 105018
rect 4330 104966 4342 105018
rect 4342 104966 4356 105018
rect 4380 104966 4394 105018
rect 4394 104966 4406 105018
rect 4406 104966 4436 105018
rect 4460 104966 4470 105018
rect 4470 104966 4516 105018
rect 4220 104964 4276 104966
rect 4300 104964 4356 104966
rect 4380 104964 4436 104966
rect 4460 104964 4516 104966
rect 4220 103930 4276 103932
rect 4300 103930 4356 103932
rect 4380 103930 4436 103932
rect 4460 103930 4516 103932
rect 4220 103878 4266 103930
rect 4266 103878 4276 103930
rect 4300 103878 4330 103930
rect 4330 103878 4342 103930
rect 4342 103878 4356 103930
rect 4380 103878 4394 103930
rect 4394 103878 4406 103930
rect 4406 103878 4436 103930
rect 4460 103878 4470 103930
rect 4470 103878 4516 103930
rect 4220 103876 4276 103878
rect 4300 103876 4356 103878
rect 4380 103876 4436 103878
rect 4460 103876 4516 103878
rect 4220 102842 4276 102844
rect 4300 102842 4356 102844
rect 4380 102842 4436 102844
rect 4460 102842 4516 102844
rect 4220 102790 4266 102842
rect 4266 102790 4276 102842
rect 4300 102790 4330 102842
rect 4330 102790 4342 102842
rect 4342 102790 4356 102842
rect 4380 102790 4394 102842
rect 4394 102790 4406 102842
rect 4406 102790 4436 102842
rect 4460 102790 4470 102842
rect 4470 102790 4516 102842
rect 4220 102788 4276 102790
rect 4300 102788 4356 102790
rect 4380 102788 4436 102790
rect 4460 102788 4516 102790
rect 4220 101754 4276 101756
rect 4300 101754 4356 101756
rect 4380 101754 4436 101756
rect 4460 101754 4516 101756
rect 4220 101702 4266 101754
rect 4266 101702 4276 101754
rect 4300 101702 4330 101754
rect 4330 101702 4342 101754
rect 4342 101702 4356 101754
rect 4380 101702 4394 101754
rect 4394 101702 4406 101754
rect 4406 101702 4436 101754
rect 4460 101702 4470 101754
rect 4470 101702 4516 101754
rect 4220 101700 4276 101702
rect 4300 101700 4356 101702
rect 4380 101700 4436 101702
rect 4460 101700 4516 101702
rect 4220 100666 4276 100668
rect 4300 100666 4356 100668
rect 4380 100666 4436 100668
rect 4460 100666 4516 100668
rect 4220 100614 4266 100666
rect 4266 100614 4276 100666
rect 4300 100614 4330 100666
rect 4330 100614 4342 100666
rect 4342 100614 4356 100666
rect 4380 100614 4394 100666
rect 4394 100614 4406 100666
rect 4406 100614 4436 100666
rect 4460 100614 4470 100666
rect 4470 100614 4516 100666
rect 4220 100612 4276 100614
rect 4300 100612 4356 100614
rect 4380 100612 4436 100614
rect 4460 100612 4516 100614
rect 4220 99578 4276 99580
rect 4300 99578 4356 99580
rect 4380 99578 4436 99580
rect 4460 99578 4516 99580
rect 4220 99526 4266 99578
rect 4266 99526 4276 99578
rect 4300 99526 4330 99578
rect 4330 99526 4342 99578
rect 4342 99526 4356 99578
rect 4380 99526 4394 99578
rect 4394 99526 4406 99578
rect 4406 99526 4436 99578
rect 4460 99526 4470 99578
rect 4470 99526 4516 99578
rect 4220 99524 4276 99526
rect 4300 99524 4356 99526
rect 4380 99524 4436 99526
rect 4460 99524 4516 99526
rect 4220 98490 4276 98492
rect 4300 98490 4356 98492
rect 4380 98490 4436 98492
rect 4460 98490 4516 98492
rect 4220 98438 4266 98490
rect 4266 98438 4276 98490
rect 4300 98438 4330 98490
rect 4330 98438 4342 98490
rect 4342 98438 4356 98490
rect 4380 98438 4394 98490
rect 4394 98438 4406 98490
rect 4406 98438 4436 98490
rect 4460 98438 4470 98490
rect 4470 98438 4516 98490
rect 4220 98436 4276 98438
rect 4300 98436 4356 98438
rect 4380 98436 4436 98438
rect 4460 98436 4516 98438
rect 4220 97402 4276 97404
rect 4300 97402 4356 97404
rect 4380 97402 4436 97404
rect 4460 97402 4516 97404
rect 4220 97350 4266 97402
rect 4266 97350 4276 97402
rect 4300 97350 4330 97402
rect 4330 97350 4342 97402
rect 4342 97350 4356 97402
rect 4380 97350 4394 97402
rect 4394 97350 4406 97402
rect 4406 97350 4436 97402
rect 4460 97350 4470 97402
rect 4470 97350 4516 97402
rect 4220 97348 4276 97350
rect 4300 97348 4356 97350
rect 4380 97348 4436 97350
rect 4460 97348 4516 97350
rect 4220 96314 4276 96316
rect 4300 96314 4356 96316
rect 4380 96314 4436 96316
rect 4460 96314 4516 96316
rect 4220 96262 4266 96314
rect 4266 96262 4276 96314
rect 4300 96262 4330 96314
rect 4330 96262 4342 96314
rect 4342 96262 4356 96314
rect 4380 96262 4394 96314
rect 4394 96262 4406 96314
rect 4406 96262 4436 96314
rect 4460 96262 4470 96314
rect 4470 96262 4516 96314
rect 4220 96260 4276 96262
rect 4300 96260 4356 96262
rect 4380 96260 4436 96262
rect 4460 96260 4516 96262
rect 4220 95226 4276 95228
rect 4300 95226 4356 95228
rect 4380 95226 4436 95228
rect 4460 95226 4516 95228
rect 4220 95174 4266 95226
rect 4266 95174 4276 95226
rect 4300 95174 4330 95226
rect 4330 95174 4342 95226
rect 4342 95174 4356 95226
rect 4380 95174 4394 95226
rect 4394 95174 4406 95226
rect 4406 95174 4436 95226
rect 4460 95174 4470 95226
rect 4470 95174 4516 95226
rect 4220 95172 4276 95174
rect 4300 95172 4356 95174
rect 4380 95172 4436 95174
rect 4460 95172 4516 95174
rect 4220 94138 4276 94140
rect 4300 94138 4356 94140
rect 4380 94138 4436 94140
rect 4460 94138 4516 94140
rect 4220 94086 4266 94138
rect 4266 94086 4276 94138
rect 4300 94086 4330 94138
rect 4330 94086 4342 94138
rect 4342 94086 4356 94138
rect 4380 94086 4394 94138
rect 4394 94086 4406 94138
rect 4406 94086 4436 94138
rect 4460 94086 4470 94138
rect 4470 94086 4516 94138
rect 4220 94084 4276 94086
rect 4300 94084 4356 94086
rect 4380 94084 4436 94086
rect 4460 94084 4516 94086
rect 4220 93050 4276 93052
rect 4300 93050 4356 93052
rect 4380 93050 4436 93052
rect 4460 93050 4516 93052
rect 4220 92998 4266 93050
rect 4266 92998 4276 93050
rect 4300 92998 4330 93050
rect 4330 92998 4342 93050
rect 4342 92998 4356 93050
rect 4380 92998 4394 93050
rect 4394 92998 4406 93050
rect 4406 92998 4436 93050
rect 4460 92998 4470 93050
rect 4470 92998 4516 93050
rect 4220 92996 4276 92998
rect 4300 92996 4356 92998
rect 4380 92996 4436 92998
rect 4460 92996 4516 92998
rect 4220 91962 4276 91964
rect 4300 91962 4356 91964
rect 4380 91962 4436 91964
rect 4460 91962 4516 91964
rect 4220 91910 4266 91962
rect 4266 91910 4276 91962
rect 4300 91910 4330 91962
rect 4330 91910 4342 91962
rect 4342 91910 4356 91962
rect 4380 91910 4394 91962
rect 4394 91910 4406 91962
rect 4406 91910 4436 91962
rect 4460 91910 4470 91962
rect 4470 91910 4516 91962
rect 4220 91908 4276 91910
rect 4300 91908 4356 91910
rect 4380 91908 4436 91910
rect 4460 91908 4516 91910
rect 4220 90874 4276 90876
rect 4300 90874 4356 90876
rect 4380 90874 4436 90876
rect 4460 90874 4516 90876
rect 4220 90822 4266 90874
rect 4266 90822 4276 90874
rect 4300 90822 4330 90874
rect 4330 90822 4342 90874
rect 4342 90822 4356 90874
rect 4380 90822 4394 90874
rect 4394 90822 4406 90874
rect 4406 90822 4436 90874
rect 4460 90822 4470 90874
rect 4470 90822 4516 90874
rect 4220 90820 4276 90822
rect 4300 90820 4356 90822
rect 4380 90820 4436 90822
rect 4460 90820 4516 90822
rect 4220 89786 4276 89788
rect 4300 89786 4356 89788
rect 4380 89786 4436 89788
rect 4460 89786 4516 89788
rect 4220 89734 4266 89786
rect 4266 89734 4276 89786
rect 4300 89734 4330 89786
rect 4330 89734 4342 89786
rect 4342 89734 4356 89786
rect 4380 89734 4394 89786
rect 4394 89734 4406 89786
rect 4406 89734 4436 89786
rect 4460 89734 4470 89786
rect 4470 89734 4516 89786
rect 4220 89732 4276 89734
rect 4300 89732 4356 89734
rect 4380 89732 4436 89734
rect 4460 89732 4516 89734
rect 4220 88698 4276 88700
rect 4300 88698 4356 88700
rect 4380 88698 4436 88700
rect 4460 88698 4516 88700
rect 4220 88646 4266 88698
rect 4266 88646 4276 88698
rect 4300 88646 4330 88698
rect 4330 88646 4342 88698
rect 4342 88646 4356 88698
rect 4380 88646 4394 88698
rect 4394 88646 4406 88698
rect 4406 88646 4436 88698
rect 4460 88646 4470 88698
rect 4470 88646 4516 88698
rect 4220 88644 4276 88646
rect 4300 88644 4356 88646
rect 4380 88644 4436 88646
rect 4460 88644 4516 88646
rect 4220 87610 4276 87612
rect 4300 87610 4356 87612
rect 4380 87610 4436 87612
rect 4460 87610 4516 87612
rect 4220 87558 4266 87610
rect 4266 87558 4276 87610
rect 4300 87558 4330 87610
rect 4330 87558 4342 87610
rect 4342 87558 4356 87610
rect 4380 87558 4394 87610
rect 4394 87558 4406 87610
rect 4406 87558 4436 87610
rect 4460 87558 4470 87610
rect 4470 87558 4516 87610
rect 4220 87556 4276 87558
rect 4300 87556 4356 87558
rect 4380 87556 4436 87558
rect 4460 87556 4516 87558
rect 4220 86522 4276 86524
rect 4300 86522 4356 86524
rect 4380 86522 4436 86524
rect 4460 86522 4516 86524
rect 4220 86470 4266 86522
rect 4266 86470 4276 86522
rect 4300 86470 4330 86522
rect 4330 86470 4342 86522
rect 4342 86470 4356 86522
rect 4380 86470 4394 86522
rect 4394 86470 4406 86522
rect 4406 86470 4436 86522
rect 4460 86470 4470 86522
rect 4470 86470 4516 86522
rect 4220 86468 4276 86470
rect 4300 86468 4356 86470
rect 4380 86468 4436 86470
rect 4460 86468 4516 86470
rect 4220 85434 4276 85436
rect 4300 85434 4356 85436
rect 4380 85434 4436 85436
rect 4460 85434 4516 85436
rect 4220 85382 4266 85434
rect 4266 85382 4276 85434
rect 4300 85382 4330 85434
rect 4330 85382 4342 85434
rect 4342 85382 4356 85434
rect 4380 85382 4394 85434
rect 4394 85382 4406 85434
rect 4406 85382 4436 85434
rect 4460 85382 4470 85434
rect 4470 85382 4516 85434
rect 4220 85380 4276 85382
rect 4300 85380 4356 85382
rect 4380 85380 4436 85382
rect 4460 85380 4516 85382
rect 4220 84346 4276 84348
rect 4300 84346 4356 84348
rect 4380 84346 4436 84348
rect 4460 84346 4516 84348
rect 4220 84294 4266 84346
rect 4266 84294 4276 84346
rect 4300 84294 4330 84346
rect 4330 84294 4342 84346
rect 4342 84294 4356 84346
rect 4380 84294 4394 84346
rect 4394 84294 4406 84346
rect 4406 84294 4436 84346
rect 4460 84294 4470 84346
rect 4470 84294 4516 84346
rect 4220 84292 4276 84294
rect 4300 84292 4356 84294
rect 4380 84292 4436 84294
rect 4460 84292 4516 84294
rect 4220 83258 4276 83260
rect 4300 83258 4356 83260
rect 4380 83258 4436 83260
rect 4460 83258 4516 83260
rect 4220 83206 4266 83258
rect 4266 83206 4276 83258
rect 4300 83206 4330 83258
rect 4330 83206 4342 83258
rect 4342 83206 4356 83258
rect 4380 83206 4394 83258
rect 4394 83206 4406 83258
rect 4406 83206 4436 83258
rect 4460 83206 4470 83258
rect 4470 83206 4516 83258
rect 4220 83204 4276 83206
rect 4300 83204 4356 83206
rect 4380 83204 4436 83206
rect 4460 83204 4516 83206
rect 4220 82170 4276 82172
rect 4300 82170 4356 82172
rect 4380 82170 4436 82172
rect 4460 82170 4516 82172
rect 4220 82118 4266 82170
rect 4266 82118 4276 82170
rect 4300 82118 4330 82170
rect 4330 82118 4342 82170
rect 4342 82118 4356 82170
rect 4380 82118 4394 82170
rect 4394 82118 4406 82170
rect 4406 82118 4436 82170
rect 4460 82118 4470 82170
rect 4470 82118 4516 82170
rect 4220 82116 4276 82118
rect 4300 82116 4356 82118
rect 4380 82116 4436 82118
rect 4460 82116 4516 82118
rect 4220 81082 4276 81084
rect 4300 81082 4356 81084
rect 4380 81082 4436 81084
rect 4460 81082 4516 81084
rect 4220 81030 4266 81082
rect 4266 81030 4276 81082
rect 4300 81030 4330 81082
rect 4330 81030 4342 81082
rect 4342 81030 4356 81082
rect 4380 81030 4394 81082
rect 4394 81030 4406 81082
rect 4406 81030 4436 81082
rect 4460 81030 4470 81082
rect 4470 81030 4516 81082
rect 4220 81028 4276 81030
rect 4300 81028 4356 81030
rect 4380 81028 4436 81030
rect 4460 81028 4516 81030
rect 4220 79994 4276 79996
rect 4300 79994 4356 79996
rect 4380 79994 4436 79996
rect 4460 79994 4516 79996
rect 4220 79942 4266 79994
rect 4266 79942 4276 79994
rect 4300 79942 4330 79994
rect 4330 79942 4342 79994
rect 4342 79942 4356 79994
rect 4380 79942 4394 79994
rect 4394 79942 4406 79994
rect 4406 79942 4436 79994
rect 4460 79942 4470 79994
rect 4470 79942 4516 79994
rect 4220 79940 4276 79942
rect 4300 79940 4356 79942
rect 4380 79940 4436 79942
rect 4460 79940 4516 79942
rect 4220 78906 4276 78908
rect 4300 78906 4356 78908
rect 4380 78906 4436 78908
rect 4460 78906 4516 78908
rect 4220 78854 4266 78906
rect 4266 78854 4276 78906
rect 4300 78854 4330 78906
rect 4330 78854 4342 78906
rect 4342 78854 4356 78906
rect 4380 78854 4394 78906
rect 4394 78854 4406 78906
rect 4406 78854 4436 78906
rect 4460 78854 4470 78906
rect 4470 78854 4516 78906
rect 4220 78852 4276 78854
rect 4300 78852 4356 78854
rect 4380 78852 4436 78854
rect 4460 78852 4516 78854
rect 1490 54476 1492 54496
rect 1492 54476 1544 54496
rect 1544 54476 1546 54496
rect 1490 54440 1546 54476
rect 1490 50360 1546 50416
rect 1582 46960 1638 47016
rect 1582 34720 1638 34776
rect 1398 31320 1454 31376
rect 1398 27240 1454 27296
rect 1398 23160 1454 23216
rect 1582 19116 1584 19136
rect 1584 19116 1636 19136
rect 1636 19116 1638 19136
rect 1582 19080 1638 19116
rect 1490 15680 1546 15736
rect 1398 11600 1454 11656
rect 1582 7520 1638 7576
rect 1858 42880 1914 42936
rect 1858 38800 1914 38856
rect 1398 3476 1400 3496
rect 1400 3476 1452 3496
rect 1452 3476 1454 3496
rect 1398 3440 1454 3476
rect 4220 77818 4276 77820
rect 4300 77818 4356 77820
rect 4380 77818 4436 77820
rect 4460 77818 4516 77820
rect 4220 77766 4266 77818
rect 4266 77766 4276 77818
rect 4300 77766 4330 77818
rect 4330 77766 4342 77818
rect 4342 77766 4356 77818
rect 4380 77766 4394 77818
rect 4394 77766 4406 77818
rect 4406 77766 4436 77818
rect 4460 77766 4470 77818
rect 4470 77766 4516 77818
rect 4220 77764 4276 77766
rect 4300 77764 4356 77766
rect 4380 77764 4436 77766
rect 4460 77764 4516 77766
rect 4220 76730 4276 76732
rect 4300 76730 4356 76732
rect 4380 76730 4436 76732
rect 4460 76730 4516 76732
rect 4220 76678 4266 76730
rect 4266 76678 4276 76730
rect 4300 76678 4330 76730
rect 4330 76678 4342 76730
rect 4342 76678 4356 76730
rect 4380 76678 4394 76730
rect 4394 76678 4406 76730
rect 4406 76678 4436 76730
rect 4460 76678 4470 76730
rect 4470 76678 4516 76730
rect 4220 76676 4276 76678
rect 4300 76676 4356 76678
rect 4380 76676 4436 76678
rect 4460 76676 4516 76678
rect 4220 75642 4276 75644
rect 4300 75642 4356 75644
rect 4380 75642 4436 75644
rect 4460 75642 4516 75644
rect 4220 75590 4266 75642
rect 4266 75590 4276 75642
rect 4300 75590 4330 75642
rect 4330 75590 4342 75642
rect 4342 75590 4356 75642
rect 4380 75590 4394 75642
rect 4394 75590 4406 75642
rect 4406 75590 4436 75642
rect 4460 75590 4470 75642
rect 4470 75590 4516 75642
rect 4220 75588 4276 75590
rect 4300 75588 4356 75590
rect 4380 75588 4436 75590
rect 4460 75588 4516 75590
rect 4220 74554 4276 74556
rect 4300 74554 4356 74556
rect 4380 74554 4436 74556
rect 4460 74554 4516 74556
rect 4220 74502 4266 74554
rect 4266 74502 4276 74554
rect 4300 74502 4330 74554
rect 4330 74502 4342 74554
rect 4342 74502 4356 74554
rect 4380 74502 4394 74554
rect 4394 74502 4406 74554
rect 4406 74502 4436 74554
rect 4460 74502 4470 74554
rect 4470 74502 4516 74554
rect 4220 74500 4276 74502
rect 4300 74500 4356 74502
rect 4380 74500 4436 74502
rect 4460 74500 4516 74502
rect 4220 73466 4276 73468
rect 4300 73466 4356 73468
rect 4380 73466 4436 73468
rect 4460 73466 4516 73468
rect 4220 73414 4266 73466
rect 4266 73414 4276 73466
rect 4300 73414 4330 73466
rect 4330 73414 4342 73466
rect 4342 73414 4356 73466
rect 4380 73414 4394 73466
rect 4394 73414 4406 73466
rect 4406 73414 4436 73466
rect 4460 73414 4470 73466
rect 4470 73414 4516 73466
rect 4220 73412 4276 73414
rect 4300 73412 4356 73414
rect 4380 73412 4436 73414
rect 4460 73412 4516 73414
rect 4220 72378 4276 72380
rect 4300 72378 4356 72380
rect 4380 72378 4436 72380
rect 4460 72378 4516 72380
rect 4220 72326 4266 72378
rect 4266 72326 4276 72378
rect 4300 72326 4330 72378
rect 4330 72326 4342 72378
rect 4342 72326 4356 72378
rect 4380 72326 4394 72378
rect 4394 72326 4406 72378
rect 4406 72326 4436 72378
rect 4460 72326 4470 72378
rect 4470 72326 4516 72378
rect 4220 72324 4276 72326
rect 4300 72324 4356 72326
rect 4380 72324 4436 72326
rect 4460 72324 4516 72326
rect 4220 71290 4276 71292
rect 4300 71290 4356 71292
rect 4380 71290 4436 71292
rect 4460 71290 4516 71292
rect 4220 71238 4266 71290
rect 4266 71238 4276 71290
rect 4300 71238 4330 71290
rect 4330 71238 4342 71290
rect 4342 71238 4356 71290
rect 4380 71238 4394 71290
rect 4394 71238 4406 71290
rect 4406 71238 4436 71290
rect 4460 71238 4470 71290
rect 4470 71238 4516 71290
rect 4220 71236 4276 71238
rect 4300 71236 4356 71238
rect 4380 71236 4436 71238
rect 4460 71236 4516 71238
rect 4220 70202 4276 70204
rect 4300 70202 4356 70204
rect 4380 70202 4436 70204
rect 4460 70202 4516 70204
rect 4220 70150 4266 70202
rect 4266 70150 4276 70202
rect 4300 70150 4330 70202
rect 4330 70150 4342 70202
rect 4342 70150 4356 70202
rect 4380 70150 4394 70202
rect 4394 70150 4406 70202
rect 4406 70150 4436 70202
rect 4460 70150 4470 70202
rect 4470 70150 4516 70202
rect 4220 70148 4276 70150
rect 4300 70148 4356 70150
rect 4380 70148 4436 70150
rect 4460 70148 4516 70150
rect 4220 69114 4276 69116
rect 4300 69114 4356 69116
rect 4380 69114 4436 69116
rect 4460 69114 4516 69116
rect 4220 69062 4266 69114
rect 4266 69062 4276 69114
rect 4300 69062 4330 69114
rect 4330 69062 4342 69114
rect 4342 69062 4356 69114
rect 4380 69062 4394 69114
rect 4394 69062 4406 69114
rect 4406 69062 4436 69114
rect 4460 69062 4470 69114
rect 4470 69062 4516 69114
rect 4220 69060 4276 69062
rect 4300 69060 4356 69062
rect 4380 69060 4436 69062
rect 4460 69060 4516 69062
rect 4220 68026 4276 68028
rect 4300 68026 4356 68028
rect 4380 68026 4436 68028
rect 4460 68026 4516 68028
rect 4220 67974 4266 68026
rect 4266 67974 4276 68026
rect 4300 67974 4330 68026
rect 4330 67974 4342 68026
rect 4342 67974 4356 68026
rect 4380 67974 4394 68026
rect 4394 67974 4406 68026
rect 4406 67974 4436 68026
rect 4460 67974 4470 68026
rect 4470 67974 4516 68026
rect 4220 67972 4276 67974
rect 4300 67972 4356 67974
rect 4380 67972 4436 67974
rect 4460 67972 4516 67974
rect 4220 66938 4276 66940
rect 4300 66938 4356 66940
rect 4380 66938 4436 66940
rect 4460 66938 4516 66940
rect 4220 66886 4266 66938
rect 4266 66886 4276 66938
rect 4300 66886 4330 66938
rect 4330 66886 4342 66938
rect 4342 66886 4356 66938
rect 4380 66886 4394 66938
rect 4394 66886 4406 66938
rect 4406 66886 4436 66938
rect 4460 66886 4470 66938
rect 4470 66886 4516 66938
rect 4220 66884 4276 66886
rect 4300 66884 4356 66886
rect 4380 66884 4436 66886
rect 4460 66884 4516 66886
rect 4220 65850 4276 65852
rect 4300 65850 4356 65852
rect 4380 65850 4436 65852
rect 4460 65850 4516 65852
rect 4220 65798 4266 65850
rect 4266 65798 4276 65850
rect 4300 65798 4330 65850
rect 4330 65798 4342 65850
rect 4342 65798 4356 65850
rect 4380 65798 4394 65850
rect 4394 65798 4406 65850
rect 4406 65798 4436 65850
rect 4460 65798 4470 65850
rect 4470 65798 4516 65850
rect 4220 65796 4276 65798
rect 4300 65796 4356 65798
rect 4380 65796 4436 65798
rect 4460 65796 4516 65798
rect 19580 117530 19636 117532
rect 19660 117530 19716 117532
rect 19740 117530 19796 117532
rect 19820 117530 19876 117532
rect 19580 117478 19626 117530
rect 19626 117478 19636 117530
rect 19660 117478 19690 117530
rect 19690 117478 19702 117530
rect 19702 117478 19716 117530
rect 19740 117478 19754 117530
rect 19754 117478 19766 117530
rect 19766 117478 19796 117530
rect 19820 117478 19830 117530
rect 19830 117478 19876 117530
rect 19580 117476 19636 117478
rect 19660 117476 19716 117478
rect 19740 117476 19796 117478
rect 19820 117476 19876 117478
rect 4220 64762 4276 64764
rect 4300 64762 4356 64764
rect 4380 64762 4436 64764
rect 4460 64762 4516 64764
rect 4220 64710 4266 64762
rect 4266 64710 4276 64762
rect 4300 64710 4330 64762
rect 4330 64710 4342 64762
rect 4342 64710 4356 64762
rect 4380 64710 4394 64762
rect 4394 64710 4406 64762
rect 4406 64710 4436 64762
rect 4460 64710 4470 64762
rect 4470 64710 4516 64762
rect 4220 64708 4276 64710
rect 4300 64708 4356 64710
rect 4380 64708 4436 64710
rect 4460 64708 4516 64710
rect 4220 63674 4276 63676
rect 4300 63674 4356 63676
rect 4380 63674 4436 63676
rect 4460 63674 4516 63676
rect 4220 63622 4266 63674
rect 4266 63622 4276 63674
rect 4300 63622 4330 63674
rect 4330 63622 4342 63674
rect 4342 63622 4356 63674
rect 4380 63622 4394 63674
rect 4394 63622 4406 63674
rect 4406 63622 4436 63674
rect 4460 63622 4470 63674
rect 4470 63622 4516 63674
rect 4220 63620 4276 63622
rect 4300 63620 4356 63622
rect 4380 63620 4436 63622
rect 4460 63620 4516 63622
rect 4220 62586 4276 62588
rect 4300 62586 4356 62588
rect 4380 62586 4436 62588
rect 4460 62586 4516 62588
rect 4220 62534 4266 62586
rect 4266 62534 4276 62586
rect 4300 62534 4330 62586
rect 4330 62534 4342 62586
rect 4342 62534 4356 62586
rect 4380 62534 4394 62586
rect 4394 62534 4406 62586
rect 4406 62534 4436 62586
rect 4460 62534 4470 62586
rect 4470 62534 4516 62586
rect 4220 62532 4276 62534
rect 4300 62532 4356 62534
rect 4380 62532 4436 62534
rect 4460 62532 4516 62534
rect 4220 61498 4276 61500
rect 4300 61498 4356 61500
rect 4380 61498 4436 61500
rect 4460 61498 4516 61500
rect 4220 61446 4266 61498
rect 4266 61446 4276 61498
rect 4300 61446 4330 61498
rect 4330 61446 4342 61498
rect 4342 61446 4356 61498
rect 4380 61446 4394 61498
rect 4394 61446 4406 61498
rect 4406 61446 4436 61498
rect 4460 61446 4470 61498
rect 4470 61446 4516 61498
rect 4220 61444 4276 61446
rect 4300 61444 4356 61446
rect 4380 61444 4436 61446
rect 4460 61444 4516 61446
rect 19580 116442 19636 116444
rect 19660 116442 19716 116444
rect 19740 116442 19796 116444
rect 19820 116442 19876 116444
rect 19580 116390 19626 116442
rect 19626 116390 19636 116442
rect 19660 116390 19690 116442
rect 19690 116390 19702 116442
rect 19702 116390 19716 116442
rect 19740 116390 19754 116442
rect 19754 116390 19766 116442
rect 19766 116390 19796 116442
rect 19820 116390 19830 116442
rect 19830 116390 19876 116442
rect 19580 116388 19636 116390
rect 19660 116388 19716 116390
rect 19740 116388 19796 116390
rect 19820 116388 19876 116390
rect 19580 115354 19636 115356
rect 19660 115354 19716 115356
rect 19740 115354 19796 115356
rect 19820 115354 19876 115356
rect 19580 115302 19626 115354
rect 19626 115302 19636 115354
rect 19660 115302 19690 115354
rect 19690 115302 19702 115354
rect 19702 115302 19716 115354
rect 19740 115302 19754 115354
rect 19754 115302 19766 115354
rect 19766 115302 19796 115354
rect 19820 115302 19830 115354
rect 19830 115302 19876 115354
rect 19580 115300 19636 115302
rect 19660 115300 19716 115302
rect 19740 115300 19796 115302
rect 19820 115300 19876 115302
rect 19580 114266 19636 114268
rect 19660 114266 19716 114268
rect 19740 114266 19796 114268
rect 19820 114266 19876 114268
rect 19580 114214 19626 114266
rect 19626 114214 19636 114266
rect 19660 114214 19690 114266
rect 19690 114214 19702 114266
rect 19702 114214 19716 114266
rect 19740 114214 19754 114266
rect 19754 114214 19766 114266
rect 19766 114214 19796 114266
rect 19820 114214 19830 114266
rect 19830 114214 19876 114266
rect 19580 114212 19636 114214
rect 19660 114212 19716 114214
rect 19740 114212 19796 114214
rect 19820 114212 19876 114214
rect 19580 113178 19636 113180
rect 19660 113178 19716 113180
rect 19740 113178 19796 113180
rect 19820 113178 19876 113180
rect 19580 113126 19626 113178
rect 19626 113126 19636 113178
rect 19660 113126 19690 113178
rect 19690 113126 19702 113178
rect 19702 113126 19716 113178
rect 19740 113126 19754 113178
rect 19754 113126 19766 113178
rect 19766 113126 19796 113178
rect 19820 113126 19830 113178
rect 19830 113126 19876 113178
rect 19580 113124 19636 113126
rect 19660 113124 19716 113126
rect 19740 113124 19796 113126
rect 19820 113124 19876 113126
rect 19580 112090 19636 112092
rect 19660 112090 19716 112092
rect 19740 112090 19796 112092
rect 19820 112090 19876 112092
rect 19580 112038 19626 112090
rect 19626 112038 19636 112090
rect 19660 112038 19690 112090
rect 19690 112038 19702 112090
rect 19702 112038 19716 112090
rect 19740 112038 19754 112090
rect 19754 112038 19766 112090
rect 19766 112038 19796 112090
rect 19820 112038 19830 112090
rect 19830 112038 19876 112090
rect 19580 112036 19636 112038
rect 19660 112036 19716 112038
rect 19740 112036 19796 112038
rect 19820 112036 19876 112038
rect 19580 111002 19636 111004
rect 19660 111002 19716 111004
rect 19740 111002 19796 111004
rect 19820 111002 19876 111004
rect 19580 110950 19626 111002
rect 19626 110950 19636 111002
rect 19660 110950 19690 111002
rect 19690 110950 19702 111002
rect 19702 110950 19716 111002
rect 19740 110950 19754 111002
rect 19754 110950 19766 111002
rect 19766 110950 19796 111002
rect 19820 110950 19830 111002
rect 19830 110950 19876 111002
rect 19580 110948 19636 110950
rect 19660 110948 19716 110950
rect 19740 110948 19796 110950
rect 19820 110948 19876 110950
rect 19580 109914 19636 109916
rect 19660 109914 19716 109916
rect 19740 109914 19796 109916
rect 19820 109914 19876 109916
rect 19580 109862 19626 109914
rect 19626 109862 19636 109914
rect 19660 109862 19690 109914
rect 19690 109862 19702 109914
rect 19702 109862 19716 109914
rect 19740 109862 19754 109914
rect 19754 109862 19766 109914
rect 19766 109862 19796 109914
rect 19820 109862 19830 109914
rect 19830 109862 19876 109914
rect 19580 109860 19636 109862
rect 19660 109860 19716 109862
rect 19740 109860 19796 109862
rect 19820 109860 19876 109862
rect 19580 108826 19636 108828
rect 19660 108826 19716 108828
rect 19740 108826 19796 108828
rect 19820 108826 19876 108828
rect 19580 108774 19626 108826
rect 19626 108774 19636 108826
rect 19660 108774 19690 108826
rect 19690 108774 19702 108826
rect 19702 108774 19716 108826
rect 19740 108774 19754 108826
rect 19754 108774 19766 108826
rect 19766 108774 19796 108826
rect 19820 108774 19830 108826
rect 19830 108774 19876 108826
rect 19580 108772 19636 108774
rect 19660 108772 19716 108774
rect 19740 108772 19796 108774
rect 19820 108772 19876 108774
rect 19580 107738 19636 107740
rect 19660 107738 19716 107740
rect 19740 107738 19796 107740
rect 19820 107738 19876 107740
rect 19580 107686 19626 107738
rect 19626 107686 19636 107738
rect 19660 107686 19690 107738
rect 19690 107686 19702 107738
rect 19702 107686 19716 107738
rect 19740 107686 19754 107738
rect 19754 107686 19766 107738
rect 19766 107686 19796 107738
rect 19820 107686 19830 107738
rect 19830 107686 19876 107738
rect 19580 107684 19636 107686
rect 19660 107684 19716 107686
rect 19740 107684 19796 107686
rect 19820 107684 19876 107686
rect 19580 106650 19636 106652
rect 19660 106650 19716 106652
rect 19740 106650 19796 106652
rect 19820 106650 19876 106652
rect 19580 106598 19626 106650
rect 19626 106598 19636 106650
rect 19660 106598 19690 106650
rect 19690 106598 19702 106650
rect 19702 106598 19716 106650
rect 19740 106598 19754 106650
rect 19754 106598 19766 106650
rect 19766 106598 19796 106650
rect 19820 106598 19830 106650
rect 19830 106598 19876 106650
rect 19580 106596 19636 106598
rect 19660 106596 19716 106598
rect 19740 106596 19796 106598
rect 19820 106596 19876 106598
rect 19580 105562 19636 105564
rect 19660 105562 19716 105564
rect 19740 105562 19796 105564
rect 19820 105562 19876 105564
rect 19580 105510 19626 105562
rect 19626 105510 19636 105562
rect 19660 105510 19690 105562
rect 19690 105510 19702 105562
rect 19702 105510 19716 105562
rect 19740 105510 19754 105562
rect 19754 105510 19766 105562
rect 19766 105510 19796 105562
rect 19820 105510 19830 105562
rect 19830 105510 19876 105562
rect 19580 105508 19636 105510
rect 19660 105508 19716 105510
rect 19740 105508 19796 105510
rect 19820 105508 19876 105510
rect 19580 104474 19636 104476
rect 19660 104474 19716 104476
rect 19740 104474 19796 104476
rect 19820 104474 19876 104476
rect 19580 104422 19626 104474
rect 19626 104422 19636 104474
rect 19660 104422 19690 104474
rect 19690 104422 19702 104474
rect 19702 104422 19716 104474
rect 19740 104422 19754 104474
rect 19754 104422 19766 104474
rect 19766 104422 19796 104474
rect 19820 104422 19830 104474
rect 19830 104422 19876 104474
rect 19580 104420 19636 104422
rect 19660 104420 19716 104422
rect 19740 104420 19796 104422
rect 19820 104420 19876 104422
rect 19580 103386 19636 103388
rect 19660 103386 19716 103388
rect 19740 103386 19796 103388
rect 19820 103386 19876 103388
rect 19580 103334 19626 103386
rect 19626 103334 19636 103386
rect 19660 103334 19690 103386
rect 19690 103334 19702 103386
rect 19702 103334 19716 103386
rect 19740 103334 19754 103386
rect 19754 103334 19766 103386
rect 19766 103334 19796 103386
rect 19820 103334 19830 103386
rect 19830 103334 19876 103386
rect 19580 103332 19636 103334
rect 19660 103332 19716 103334
rect 19740 103332 19796 103334
rect 19820 103332 19876 103334
rect 19580 102298 19636 102300
rect 19660 102298 19716 102300
rect 19740 102298 19796 102300
rect 19820 102298 19876 102300
rect 19580 102246 19626 102298
rect 19626 102246 19636 102298
rect 19660 102246 19690 102298
rect 19690 102246 19702 102298
rect 19702 102246 19716 102298
rect 19740 102246 19754 102298
rect 19754 102246 19766 102298
rect 19766 102246 19796 102298
rect 19820 102246 19830 102298
rect 19830 102246 19876 102298
rect 19580 102244 19636 102246
rect 19660 102244 19716 102246
rect 19740 102244 19796 102246
rect 19820 102244 19876 102246
rect 19580 101210 19636 101212
rect 19660 101210 19716 101212
rect 19740 101210 19796 101212
rect 19820 101210 19876 101212
rect 19580 101158 19626 101210
rect 19626 101158 19636 101210
rect 19660 101158 19690 101210
rect 19690 101158 19702 101210
rect 19702 101158 19716 101210
rect 19740 101158 19754 101210
rect 19754 101158 19766 101210
rect 19766 101158 19796 101210
rect 19820 101158 19830 101210
rect 19830 101158 19876 101210
rect 19580 101156 19636 101158
rect 19660 101156 19716 101158
rect 19740 101156 19796 101158
rect 19820 101156 19876 101158
rect 19580 100122 19636 100124
rect 19660 100122 19716 100124
rect 19740 100122 19796 100124
rect 19820 100122 19876 100124
rect 19580 100070 19626 100122
rect 19626 100070 19636 100122
rect 19660 100070 19690 100122
rect 19690 100070 19702 100122
rect 19702 100070 19716 100122
rect 19740 100070 19754 100122
rect 19754 100070 19766 100122
rect 19766 100070 19796 100122
rect 19820 100070 19830 100122
rect 19830 100070 19876 100122
rect 19580 100068 19636 100070
rect 19660 100068 19716 100070
rect 19740 100068 19796 100070
rect 19820 100068 19876 100070
rect 19580 99034 19636 99036
rect 19660 99034 19716 99036
rect 19740 99034 19796 99036
rect 19820 99034 19876 99036
rect 19580 98982 19626 99034
rect 19626 98982 19636 99034
rect 19660 98982 19690 99034
rect 19690 98982 19702 99034
rect 19702 98982 19716 99034
rect 19740 98982 19754 99034
rect 19754 98982 19766 99034
rect 19766 98982 19796 99034
rect 19820 98982 19830 99034
rect 19830 98982 19876 99034
rect 19580 98980 19636 98982
rect 19660 98980 19716 98982
rect 19740 98980 19796 98982
rect 19820 98980 19876 98982
rect 19580 97946 19636 97948
rect 19660 97946 19716 97948
rect 19740 97946 19796 97948
rect 19820 97946 19876 97948
rect 19580 97894 19626 97946
rect 19626 97894 19636 97946
rect 19660 97894 19690 97946
rect 19690 97894 19702 97946
rect 19702 97894 19716 97946
rect 19740 97894 19754 97946
rect 19754 97894 19766 97946
rect 19766 97894 19796 97946
rect 19820 97894 19830 97946
rect 19830 97894 19876 97946
rect 19580 97892 19636 97894
rect 19660 97892 19716 97894
rect 19740 97892 19796 97894
rect 19820 97892 19876 97894
rect 19580 96858 19636 96860
rect 19660 96858 19716 96860
rect 19740 96858 19796 96860
rect 19820 96858 19876 96860
rect 19580 96806 19626 96858
rect 19626 96806 19636 96858
rect 19660 96806 19690 96858
rect 19690 96806 19702 96858
rect 19702 96806 19716 96858
rect 19740 96806 19754 96858
rect 19754 96806 19766 96858
rect 19766 96806 19796 96858
rect 19820 96806 19830 96858
rect 19830 96806 19876 96858
rect 19580 96804 19636 96806
rect 19660 96804 19716 96806
rect 19740 96804 19796 96806
rect 19820 96804 19876 96806
rect 19580 95770 19636 95772
rect 19660 95770 19716 95772
rect 19740 95770 19796 95772
rect 19820 95770 19876 95772
rect 19580 95718 19626 95770
rect 19626 95718 19636 95770
rect 19660 95718 19690 95770
rect 19690 95718 19702 95770
rect 19702 95718 19716 95770
rect 19740 95718 19754 95770
rect 19754 95718 19766 95770
rect 19766 95718 19796 95770
rect 19820 95718 19830 95770
rect 19830 95718 19876 95770
rect 19580 95716 19636 95718
rect 19660 95716 19716 95718
rect 19740 95716 19796 95718
rect 19820 95716 19876 95718
rect 19580 94682 19636 94684
rect 19660 94682 19716 94684
rect 19740 94682 19796 94684
rect 19820 94682 19876 94684
rect 19580 94630 19626 94682
rect 19626 94630 19636 94682
rect 19660 94630 19690 94682
rect 19690 94630 19702 94682
rect 19702 94630 19716 94682
rect 19740 94630 19754 94682
rect 19754 94630 19766 94682
rect 19766 94630 19796 94682
rect 19820 94630 19830 94682
rect 19830 94630 19876 94682
rect 19580 94628 19636 94630
rect 19660 94628 19716 94630
rect 19740 94628 19796 94630
rect 19820 94628 19876 94630
rect 19580 93594 19636 93596
rect 19660 93594 19716 93596
rect 19740 93594 19796 93596
rect 19820 93594 19876 93596
rect 19580 93542 19626 93594
rect 19626 93542 19636 93594
rect 19660 93542 19690 93594
rect 19690 93542 19702 93594
rect 19702 93542 19716 93594
rect 19740 93542 19754 93594
rect 19754 93542 19766 93594
rect 19766 93542 19796 93594
rect 19820 93542 19830 93594
rect 19830 93542 19876 93594
rect 19580 93540 19636 93542
rect 19660 93540 19716 93542
rect 19740 93540 19796 93542
rect 19820 93540 19876 93542
rect 19580 92506 19636 92508
rect 19660 92506 19716 92508
rect 19740 92506 19796 92508
rect 19820 92506 19876 92508
rect 19580 92454 19626 92506
rect 19626 92454 19636 92506
rect 19660 92454 19690 92506
rect 19690 92454 19702 92506
rect 19702 92454 19716 92506
rect 19740 92454 19754 92506
rect 19754 92454 19766 92506
rect 19766 92454 19796 92506
rect 19820 92454 19830 92506
rect 19830 92454 19876 92506
rect 19580 92452 19636 92454
rect 19660 92452 19716 92454
rect 19740 92452 19796 92454
rect 19820 92452 19876 92454
rect 19580 91418 19636 91420
rect 19660 91418 19716 91420
rect 19740 91418 19796 91420
rect 19820 91418 19876 91420
rect 19580 91366 19626 91418
rect 19626 91366 19636 91418
rect 19660 91366 19690 91418
rect 19690 91366 19702 91418
rect 19702 91366 19716 91418
rect 19740 91366 19754 91418
rect 19754 91366 19766 91418
rect 19766 91366 19796 91418
rect 19820 91366 19830 91418
rect 19830 91366 19876 91418
rect 19580 91364 19636 91366
rect 19660 91364 19716 91366
rect 19740 91364 19796 91366
rect 19820 91364 19876 91366
rect 19580 90330 19636 90332
rect 19660 90330 19716 90332
rect 19740 90330 19796 90332
rect 19820 90330 19876 90332
rect 19580 90278 19626 90330
rect 19626 90278 19636 90330
rect 19660 90278 19690 90330
rect 19690 90278 19702 90330
rect 19702 90278 19716 90330
rect 19740 90278 19754 90330
rect 19754 90278 19766 90330
rect 19766 90278 19796 90330
rect 19820 90278 19830 90330
rect 19830 90278 19876 90330
rect 19580 90276 19636 90278
rect 19660 90276 19716 90278
rect 19740 90276 19796 90278
rect 19820 90276 19876 90278
rect 19580 89242 19636 89244
rect 19660 89242 19716 89244
rect 19740 89242 19796 89244
rect 19820 89242 19876 89244
rect 19580 89190 19626 89242
rect 19626 89190 19636 89242
rect 19660 89190 19690 89242
rect 19690 89190 19702 89242
rect 19702 89190 19716 89242
rect 19740 89190 19754 89242
rect 19754 89190 19766 89242
rect 19766 89190 19796 89242
rect 19820 89190 19830 89242
rect 19830 89190 19876 89242
rect 19580 89188 19636 89190
rect 19660 89188 19716 89190
rect 19740 89188 19796 89190
rect 19820 89188 19876 89190
rect 19580 88154 19636 88156
rect 19660 88154 19716 88156
rect 19740 88154 19796 88156
rect 19820 88154 19876 88156
rect 19580 88102 19626 88154
rect 19626 88102 19636 88154
rect 19660 88102 19690 88154
rect 19690 88102 19702 88154
rect 19702 88102 19716 88154
rect 19740 88102 19754 88154
rect 19754 88102 19766 88154
rect 19766 88102 19796 88154
rect 19820 88102 19830 88154
rect 19830 88102 19876 88154
rect 19580 88100 19636 88102
rect 19660 88100 19716 88102
rect 19740 88100 19796 88102
rect 19820 88100 19876 88102
rect 19580 87066 19636 87068
rect 19660 87066 19716 87068
rect 19740 87066 19796 87068
rect 19820 87066 19876 87068
rect 19580 87014 19626 87066
rect 19626 87014 19636 87066
rect 19660 87014 19690 87066
rect 19690 87014 19702 87066
rect 19702 87014 19716 87066
rect 19740 87014 19754 87066
rect 19754 87014 19766 87066
rect 19766 87014 19796 87066
rect 19820 87014 19830 87066
rect 19830 87014 19876 87066
rect 19580 87012 19636 87014
rect 19660 87012 19716 87014
rect 19740 87012 19796 87014
rect 19820 87012 19876 87014
rect 19580 85978 19636 85980
rect 19660 85978 19716 85980
rect 19740 85978 19796 85980
rect 19820 85978 19876 85980
rect 19580 85926 19626 85978
rect 19626 85926 19636 85978
rect 19660 85926 19690 85978
rect 19690 85926 19702 85978
rect 19702 85926 19716 85978
rect 19740 85926 19754 85978
rect 19754 85926 19766 85978
rect 19766 85926 19796 85978
rect 19820 85926 19830 85978
rect 19830 85926 19876 85978
rect 19580 85924 19636 85926
rect 19660 85924 19716 85926
rect 19740 85924 19796 85926
rect 19820 85924 19876 85926
rect 19580 84890 19636 84892
rect 19660 84890 19716 84892
rect 19740 84890 19796 84892
rect 19820 84890 19876 84892
rect 19580 84838 19626 84890
rect 19626 84838 19636 84890
rect 19660 84838 19690 84890
rect 19690 84838 19702 84890
rect 19702 84838 19716 84890
rect 19740 84838 19754 84890
rect 19754 84838 19766 84890
rect 19766 84838 19796 84890
rect 19820 84838 19830 84890
rect 19830 84838 19876 84890
rect 19580 84836 19636 84838
rect 19660 84836 19716 84838
rect 19740 84836 19796 84838
rect 19820 84836 19876 84838
rect 19580 83802 19636 83804
rect 19660 83802 19716 83804
rect 19740 83802 19796 83804
rect 19820 83802 19876 83804
rect 19580 83750 19626 83802
rect 19626 83750 19636 83802
rect 19660 83750 19690 83802
rect 19690 83750 19702 83802
rect 19702 83750 19716 83802
rect 19740 83750 19754 83802
rect 19754 83750 19766 83802
rect 19766 83750 19796 83802
rect 19820 83750 19830 83802
rect 19830 83750 19876 83802
rect 19580 83748 19636 83750
rect 19660 83748 19716 83750
rect 19740 83748 19796 83750
rect 19820 83748 19876 83750
rect 19580 82714 19636 82716
rect 19660 82714 19716 82716
rect 19740 82714 19796 82716
rect 19820 82714 19876 82716
rect 19580 82662 19626 82714
rect 19626 82662 19636 82714
rect 19660 82662 19690 82714
rect 19690 82662 19702 82714
rect 19702 82662 19716 82714
rect 19740 82662 19754 82714
rect 19754 82662 19766 82714
rect 19766 82662 19796 82714
rect 19820 82662 19830 82714
rect 19830 82662 19876 82714
rect 19580 82660 19636 82662
rect 19660 82660 19716 82662
rect 19740 82660 19796 82662
rect 19820 82660 19876 82662
rect 19580 81626 19636 81628
rect 19660 81626 19716 81628
rect 19740 81626 19796 81628
rect 19820 81626 19876 81628
rect 19580 81574 19626 81626
rect 19626 81574 19636 81626
rect 19660 81574 19690 81626
rect 19690 81574 19702 81626
rect 19702 81574 19716 81626
rect 19740 81574 19754 81626
rect 19754 81574 19766 81626
rect 19766 81574 19796 81626
rect 19820 81574 19830 81626
rect 19830 81574 19876 81626
rect 19580 81572 19636 81574
rect 19660 81572 19716 81574
rect 19740 81572 19796 81574
rect 19820 81572 19876 81574
rect 19580 80538 19636 80540
rect 19660 80538 19716 80540
rect 19740 80538 19796 80540
rect 19820 80538 19876 80540
rect 19580 80486 19626 80538
rect 19626 80486 19636 80538
rect 19660 80486 19690 80538
rect 19690 80486 19702 80538
rect 19702 80486 19716 80538
rect 19740 80486 19754 80538
rect 19754 80486 19766 80538
rect 19766 80486 19796 80538
rect 19820 80486 19830 80538
rect 19830 80486 19876 80538
rect 19580 80484 19636 80486
rect 19660 80484 19716 80486
rect 19740 80484 19796 80486
rect 19820 80484 19876 80486
rect 19580 79450 19636 79452
rect 19660 79450 19716 79452
rect 19740 79450 19796 79452
rect 19820 79450 19876 79452
rect 19580 79398 19626 79450
rect 19626 79398 19636 79450
rect 19660 79398 19690 79450
rect 19690 79398 19702 79450
rect 19702 79398 19716 79450
rect 19740 79398 19754 79450
rect 19754 79398 19766 79450
rect 19766 79398 19796 79450
rect 19820 79398 19830 79450
rect 19830 79398 19876 79450
rect 19580 79396 19636 79398
rect 19660 79396 19716 79398
rect 19740 79396 19796 79398
rect 19820 79396 19876 79398
rect 19580 78362 19636 78364
rect 19660 78362 19716 78364
rect 19740 78362 19796 78364
rect 19820 78362 19876 78364
rect 19580 78310 19626 78362
rect 19626 78310 19636 78362
rect 19660 78310 19690 78362
rect 19690 78310 19702 78362
rect 19702 78310 19716 78362
rect 19740 78310 19754 78362
rect 19754 78310 19766 78362
rect 19766 78310 19796 78362
rect 19820 78310 19830 78362
rect 19830 78310 19876 78362
rect 19580 78308 19636 78310
rect 19660 78308 19716 78310
rect 19740 78308 19796 78310
rect 19820 78308 19876 78310
rect 19580 77274 19636 77276
rect 19660 77274 19716 77276
rect 19740 77274 19796 77276
rect 19820 77274 19876 77276
rect 19580 77222 19626 77274
rect 19626 77222 19636 77274
rect 19660 77222 19690 77274
rect 19690 77222 19702 77274
rect 19702 77222 19716 77274
rect 19740 77222 19754 77274
rect 19754 77222 19766 77274
rect 19766 77222 19796 77274
rect 19820 77222 19830 77274
rect 19830 77222 19876 77274
rect 19580 77220 19636 77222
rect 19660 77220 19716 77222
rect 19740 77220 19796 77222
rect 19820 77220 19876 77222
rect 19580 76186 19636 76188
rect 19660 76186 19716 76188
rect 19740 76186 19796 76188
rect 19820 76186 19876 76188
rect 19580 76134 19626 76186
rect 19626 76134 19636 76186
rect 19660 76134 19690 76186
rect 19690 76134 19702 76186
rect 19702 76134 19716 76186
rect 19740 76134 19754 76186
rect 19754 76134 19766 76186
rect 19766 76134 19796 76186
rect 19820 76134 19830 76186
rect 19830 76134 19876 76186
rect 19580 76132 19636 76134
rect 19660 76132 19716 76134
rect 19740 76132 19796 76134
rect 19820 76132 19876 76134
rect 19580 75098 19636 75100
rect 19660 75098 19716 75100
rect 19740 75098 19796 75100
rect 19820 75098 19876 75100
rect 19580 75046 19626 75098
rect 19626 75046 19636 75098
rect 19660 75046 19690 75098
rect 19690 75046 19702 75098
rect 19702 75046 19716 75098
rect 19740 75046 19754 75098
rect 19754 75046 19766 75098
rect 19766 75046 19796 75098
rect 19820 75046 19830 75098
rect 19830 75046 19876 75098
rect 19580 75044 19636 75046
rect 19660 75044 19716 75046
rect 19740 75044 19796 75046
rect 19820 75044 19876 75046
rect 19580 74010 19636 74012
rect 19660 74010 19716 74012
rect 19740 74010 19796 74012
rect 19820 74010 19876 74012
rect 19580 73958 19626 74010
rect 19626 73958 19636 74010
rect 19660 73958 19690 74010
rect 19690 73958 19702 74010
rect 19702 73958 19716 74010
rect 19740 73958 19754 74010
rect 19754 73958 19766 74010
rect 19766 73958 19796 74010
rect 19820 73958 19830 74010
rect 19830 73958 19876 74010
rect 19580 73956 19636 73958
rect 19660 73956 19716 73958
rect 19740 73956 19796 73958
rect 19820 73956 19876 73958
rect 19580 72922 19636 72924
rect 19660 72922 19716 72924
rect 19740 72922 19796 72924
rect 19820 72922 19876 72924
rect 19580 72870 19626 72922
rect 19626 72870 19636 72922
rect 19660 72870 19690 72922
rect 19690 72870 19702 72922
rect 19702 72870 19716 72922
rect 19740 72870 19754 72922
rect 19754 72870 19766 72922
rect 19766 72870 19796 72922
rect 19820 72870 19830 72922
rect 19830 72870 19876 72922
rect 19580 72868 19636 72870
rect 19660 72868 19716 72870
rect 19740 72868 19796 72870
rect 19820 72868 19876 72870
rect 19580 71834 19636 71836
rect 19660 71834 19716 71836
rect 19740 71834 19796 71836
rect 19820 71834 19876 71836
rect 19580 71782 19626 71834
rect 19626 71782 19636 71834
rect 19660 71782 19690 71834
rect 19690 71782 19702 71834
rect 19702 71782 19716 71834
rect 19740 71782 19754 71834
rect 19754 71782 19766 71834
rect 19766 71782 19796 71834
rect 19820 71782 19830 71834
rect 19830 71782 19876 71834
rect 19580 71780 19636 71782
rect 19660 71780 19716 71782
rect 19740 71780 19796 71782
rect 19820 71780 19876 71782
rect 19580 70746 19636 70748
rect 19660 70746 19716 70748
rect 19740 70746 19796 70748
rect 19820 70746 19876 70748
rect 19580 70694 19626 70746
rect 19626 70694 19636 70746
rect 19660 70694 19690 70746
rect 19690 70694 19702 70746
rect 19702 70694 19716 70746
rect 19740 70694 19754 70746
rect 19754 70694 19766 70746
rect 19766 70694 19796 70746
rect 19820 70694 19830 70746
rect 19830 70694 19876 70746
rect 19580 70692 19636 70694
rect 19660 70692 19716 70694
rect 19740 70692 19796 70694
rect 19820 70692 19876 70694
rect 19580 69658 19636 69660
rect 19660 69658 19716 69660
rect 19740 69658 19796 69660
rect 19820 69658 19876 69660
rect 19580 69606 19626 69658
rect 19626 69606 19636 69658
rect 19660 69606 19690 69658
rect 19690 69606 19702 69658
rect 19702 69606 19716 69658
rect 19740 69606 19754 69658
rect 19754 69606 19766 69658
rect 19766 69606 19796 69658
rect 19820 69606 19830 69658
rect 19830 69606 19876 69658
rect 19580 69604 19636 69606
rect 19660 69604 19716 69606
rect 19740 69604 19796 69606
rect 19820 69604 19876 69606
rect 19580 68570 19636 68572
rect 19660 68570 19716 68572
rect 19740 68570 19796 68572
rect 19820 68570 19876 68572
rect 19580 68518 19626 68570
rect 19626 68518 19636 68570
rect 19660 68518 19690 68570
rect 19690 68518 19702 68570
rect 19702 68518 19716 68570
rect 19740 68518 19754 68570
rect 19754 68518 19766 68570
rect 19766 68518 19796 68570
rect 19820 68518 19830 68570
rect 19830 68518 19876 68570
rect 19580 68516 19636 68518
rect 19660 68516 19716 68518
rect 19740 68516 19796 68518
rect 19820 68516 19876 68518
rect 19580 67482 19636 67484
rect 19660 67482 19716 67484
rect 19740 67482 19796 67484
rect 19820 67482 19876 67484
rect 19580 67430 19626 67482
rect 19626 67430 19636 67482
rect 19660 67430 19690 67482
rect 19690 67430 19702 67482
rect 19702 67430 19716 67482
rect 19740 67430 19754 67482
rect 19754 67430 19766 67482
rect 19766 67430 19796 67482
rect 19820 67430 19830 67482
rect 19830 67430 19876 67482
rect 19580 67428 19636 67430
rect 19660 67428 19716 67430
rect 19740 67428 19796 67430
rect 19820 67428 19876 67430
rect 19580 66394 19636 66396
rect 19660 66394 19716 66396
rect 19740 66394 19796 66396
rect 19820 66394 19876 66396
rect 19580 66342 19626 66394
rect 19626 66342 19636 66394
rect 19660 66342 19690 66394
rect 19690 66342 19702 66394
rect 19702 66342 19716 66394
rect 19740 66342 19754 66394
rect 19754 66342 19766 66394
rect 19766 66342 19796 66394
rect 19820 66342 19830 66394
rect 19830 66342 19876 66394
rect 19580 66340 19636 66342
rect 19660 66340 19716 66342
rect 19740 66340 19796 66342
rect 19820 66340 19876 66342
rect 19580 65306 19636 65308
rect 19660 65306 19716 65308
rect 19740 65306 19796 65308
rect 19820 65306 19876 65308
rect 19580 65254 19626 65306
rect 19626 65254 19636 65306
rect 19660 65254 19690 65306
rect 19690 65254 19702 65306
rect 19702 65254 19716 65306
rect 19740 65254 19754 65306
rect 19754 65254 19766 65306
rect 19766 65254 19796 65306
rect 19820 65254 19830 65306
rect 19830 65254 19876 65306
rect 19580 65252 19636 65254
rect 19660 65252 19716 65254
rect 19740 65252 19796 65254
rect 19820 65252 19876 65254
rect 19580 64218 19636 64220
rect 19660 64218 19716 64220
rect 19740 64218 19796 64220
rect 19820 64218 19876 64220
rect 19580 64166 19626 64218
rect 19626 64166 19636 64218
rect 19660 64166 19690 64218
rect 19690 64166 19702 64218
rect 19702 64166 19716 64218
rect 19740 64166 19754 64218
rect 19754 64166 19766 64218
rect 19766 64166 19796 64218
rect 19820 64166 19830 64218
rect 19830 64166 19876 64218
rect 19580 64164 19636 64166
rect 19660 64164 19716 64166
rect 19740 64164 19796 64166
rect 19820 64164 19876 64166
rect 19580 63130 19636 63132
rect 19660 63130 19716 63132
rect 19740 63130 19796 63132
rect 19820 63130 19876 63132
rect 19580 63078 19626 63130
rect 19626 63078 19636 63130
rect 19660 63078 19690 63130
rect 19690 63078 19702 63130
rect 19702 63078 19716 63130
rect 19740 63078 19754 63130
rect 19754 63078 19766 63130
rect 19766 63078 19796 63130
rect 19820 63078 19830 63130
rect 19830 63078 19876 63130
rect 19580 63076 19636 63078
rect 19660 63076 19716 63078
rect 19740 63076 19796 63078
rect 19820 63076 19876 63078
rect 19580 62042 19636 62044
rect 19660 62042 19716 62044
rect 19740 62042 19796 62044
rect 19820 62042 19876 62044
rect 19580 61990 19626 62042
rect 19626 61990 19636 62042
rect 19660 61990 19690 62042
rect 19690 61990 19702 62042
rect 19702 61990 19716 62042
rect 19740 61990 19754 62042
rect 19754 61990 19766 62042
rect 19766 61990 19796 62042
rect 19820 61990 19830 62042
rect 19830 61990 19876 62042
rect 19580 61988 19636 61990
rect 19660 61988 19716 61990
rect 19740 61988 19796 61990
rect 19820 61988 19876 61990
rect 19580 60954 19636 60956
rect 19660 60954 19716 60956
rect 19740 60954 19796 60956
rect 19820 60954 19876 60956
rect 19580 60902 19626 60954
rect 19626 60902 19636 60954
rect 19660 60902 19690 60954
rect 19690 60902 19702 60954
rect 19702 60902 19716 60954
rect 19740 60902 19754 60954
rect 19754 60902 19766 60954
rect 19766 60902 19796 60954
rect 19820 60902 19830 60954
rect 19830 60902 19876 60954
rect 19580 60900 19636 60902
rect 19660 60900 19716 60902
rect 19740 60900 19796 60902
rect 19820 60900 19876 60902
rect 4220 60410 4276 60412
rect 4300 60410 4356 60412
rect 4380 60410 4436 60412
rect 4460 60410 4516 60412
rect 4220 60358 4266 60410
rect 4266 60358 4276 60410
rect 4300 60358 4330 60410
rect 4330 60358 4342 60410
rect 4342 60358 4356 60410
rect 4380 60358 4394 60410
rect 4394 60358 4406 60410
rect 4406 60358 4436 60410
rect 4460 60358 4470 60410
rect 4470 60358 4516 60410
rect 4220 60356 4276 60358
rect 4300 60356 4356 60358
rect 4380 60356 4436 60358
rect 4460 60356 4516 60358
rect 34940 116986 34996 116988
rect 35020 116986 35076 116988
rect 35100 116986 35156 116988
rect 35180 116986 35236 116988
rect 34940 116934 34986 116986
rect 34986 116934 34996 116986
rect 35020 116934 35050 116986
rect 35050 116934 35062 116986
rect 35062 116934 35076 116986
rect 35100 116934 35114 116986
rect 35114 116934 35126 116986
rect 35126 116934 35156 116986
rect 35180 116934 35190 116986
rect 35190 116934 35236 116986
rect 34940 116932 34996 116934
rect 35020 116932 35076 116934
rect 35100 116932 35156 116934
rect 35180 116932 35236 116934
rect 34940 115898 34996 115900
rect 35020 115898 35076 115900
rect 35100 115898 35156 115900
rect 35180 115898 35236 115900
rect 34940 115846 34986 115898
rect 34986 115846 34996 115898
rect 35020 115846 35050 115898
rect 35050 115846 35062 115898
rect 35062 115846 35076 115898
rect 35100 115846 35114 115898
rect 35114 115846 35126 115898
rect 35126 115846 35156 115898
rect 35180 115846 35190 115898
rect 35190 115846 35236 115898
rect 34940 115844 34996 115846
rect 35020 115844 35076 115846
rect 35100 115844 35156 115846
rect 35180 115844 35236 115846
rect 34940 114810 34996 114812
rect 35020 114810 35076 114812
rect 35100 114810 35156 114812
rect 35180 114810 35236 114812
rect 34940 114758 34986 114810
rect 34986 114758 34996 114810
rect 35020 114758 35050 114810
rect 35050 114758 35062 114810
rect 35062 114758 35076 114810
rect 35100 114758 35114 114810
rect 35114 114758 35126 114810
rect 35126 114758 35156 114810
rect 35180 114758 35190 114810
rect 35190 114758 35236 114810
rect 34940 114756 34996 114758
rect 35020 114756 35076 114758
rect 35100 114756 35156 114758
rect 35180 114756 35236 114758
rect 34940 113722 34996 113724
rect 35020 113722 35076 113724
rect 35100 113722 35156 113724
rect 35180 113722 35236 113724
rect 34940 113670 34986 113722
rect 34986 113670 34996 113722
rect 35020 113670 35050 113722
rect 35050 113670 35062 113722
rect 35062 113670 35076 113722
rect 35100 113670 35114 113722
rect 35114 113670 35126 113722
rect 35126 113670 35156 113722
rect 35180 113670 35190 113722
rect 35190 113670 35236 113722
rect 34940 113668 34996 113670
rect 35020 113668 35076 113670
rect 35100 113668 35156 113670
rect 35180 113668 35236 113670
rect 34940 112634 34996 112636
rect 35020 112634 35076 112636
rect 35100 112634 35156 112636
rect 35180 112634 35236 112636
rect 34940 112582 34986 112634
rect 34986 112582 34996 112634
rect 35020 112582 35050 112634
rect 35050 112582 35062 112634
rect 35062 112582 35076 112634
rect 35100 112582 35114 112634
rect 35114 112582 35126 112634
rect 35126 112582 35156 112634
rect 35180 112582 35190 112634
rect 35190 112582 35236 112634
rect 34940 112580 34996 112582
rect 35020 112580 35076 112582
rect 35100 112580 35156 112582
rect 35180 112580 35236 112582
rect 34940 111546 34996 111548
rect 35020 111546 35076 111548
rect 35100 111546 35156 111548
rect 35180 111546 35236 111548
rect 34940 111494 34986 111546
rect 34986 111494 34996 111546
rect 35020 111494 35050 111546
rect 35050 111494 35062 111546
rect 35062 111494 35076 111546
rect 35100 111494 35114 111546
rect 35114 111494 35126 111546
rect 35126 111494 35156 111546
rect 35180 111494 35190 111546
rect 35190 111494 35236 111546
rect 34940 111492 34996 111494
rect 35020 111492 35076 111494
rect 35100 111492 35156 111494
rect 35180 111492 35236 111494
rect 34940 110458 34996 110460
rect 35020 110458 35076 110460
rect 35100 110458 35156 110460
rect 35180 110458 35236 110460
rect 34940 110406 34986 110458
rect 34986 110406 34996 110458
rect 35020 110406 35050 110458
rect 35050 110406 35062 110458
rect 35062 110406 35076 110458
rect 35100 110406 35114 110458
rect 35114 110406 35126 110458
rect 35126 110406 35156 110458
rect 35180 110406 35190 110458
rect 35190 110406 35236 110458
rect 34940 110404 34996 110406
rect 35020 110404 35076 110406
rect 35100 110404 35156 110406
rect 35180 110404 35236 110406
rect 34940 109370 34996 109372
rect 35020 109370 35076 109372
rect 35100 109370 35156 109372
rect 35180 109370 35236 109372
rect 34940 109318 34986 109370
rect 34986 109318 34996 109370
rect 35020 109318 35050 109370
rect 35050 109318 35062 109370
rect 35062 109318 35076 109370
rect 35100 109318 35114 109370
rect 35114 109318 35126 109370
rect 35126 109318 35156 109370
rect 35180 109318 35190 109370
rect 35190 109318 35236 109370
rect 34940 109316 34996 109318
rect 35020 109316 35076 109318
rect 35100 109316 35156 109318
rect 35180 109316 35236 109318
rect 34940 108282 34996 108284
rect 35020 108282 35076 108284
rect 35100 108282 35156 108284
rect 35180 108282 35236 108284
rect 34940 108230 34986 108282
rect 34986 108230 34996 108282
rect 35020 108230 35050 108282
rect 35050 108230 35062 108282
rect 35062 108230 35076 108282
rect 35100 108230 35114 108282
rect 35114 108230 35126 108282
rect 35126 108230 35156 108282
rect 35180 108230 35190 108282
rect 35190 108230 35236 108282
rect 34940 108228 34996 108230
rect 35020 108228 35076 108230
rect 35100 108228 35156 108230
rect 35180 108228 35236 108230
rect 34940 107194 34996 107196
rect 35020 107194 35076 107196
rect 35100 107194 35156 107196
rect 35180 107194 35236 107196
rect 34940 107142 34986 107194
rect 34986 107142 34996 107194
rect 35020 107142 35050 107194
rect 35050 107142 35062 107194
rect 35062 107142 35076 107194
rect 35100 107142 35114 107194
rect 35114 107142 35126 107194
rect 35126 107142 35156 107194
rect 35180 107142 35190 107194
rect 35190 107142 35236 107194
rect 34940 107140 34996 107142
rect 35020 107140 35076 107142
rect 35100 107140 35156 107142
rect 35180 107140 35236 107142
rect 34940 106106 34996 106108
rect 35020 106106 35076 106108
rect 35100 106106 35156 106108
rect 35180 106106 35236 106108
rect 34940 106054 34986 106106
rect 34986 106054 34996 106106
rect 35020 106054 35050 106106
rect 35050 106054 35062 106106
rect 35062 106054 35076 106106
rect 35100 106054 35114 106106
rect 35114 106054 35126 106106
rect 35126 106054 35156 106106
rect 35180 106054 35190 106106
rect 35190 106054 35236 106106
rect 34940 106052 34996 106054
rect 35020 106052 35076 106054
rect 35100 106052 35156 106054
rect 35180 106052 35236 106054
rect 34940 105018 34996 105020
rect 35020 105018 35076 105020
rect 35100 105018 35156 105020
rect 35180 105018 35236 105020
rect 34940 104966 34986 105018
rect 34986 104966 34996 105018
rect 35020 104966 35050 105018
rect 35050 104966 35062 105018
rect 35062 104966 35076 105018
rect 35100 104966 35114 105018
rect 35114 104966 35126 105018
rect 35126 104966 35156 105018
rect 35180 104966 35190 105018
rect 35190 104966 35236 105018
rect 34940 104964 34996 104966
rect 35020 104964 35076 104966
rect 35100 104964 35156 104966
rect 35180 104964 35236 104966
rect 34940 103930 34996 103932
rect 35020 103930 35076 103932
rect 35100 103930 35156 103932
rect 35180 103930 35236 103932
rect 34940 103878 34986 103930
rect 34986 103878 34996 103930
rect 35020 103878 35050 103930
rect 35050 103878 35062 103930
rect 35062 103878 35076 103930
rect 35100 103878 35114 103930
rect 35114 103878 35126 103930
rect 35126 103878 35156 103930
rect 35180 103878 35190 103930
rect 35190 103878 35236 103930
rect 34940 103876 34996 103878
rect 35020 103876 35076 103878
rect 35100 103876 35156 103878
rect 35180 103876 35236 103878
rect 34940 102842 34996 102844
rect 35020 102842 35076 102844
rect 35100 102842 35156 102844
rect 35180 102842 35236 102844
rect 34940 102790 34986 102842
rect 34986 102790 34996 102842
rect 35020 102790 35050 102842
rect 35050 102790 35062 102842
rect 35062 102790 35076 102842
rect 35100 102790 35114 102842
rect 35114 102790 35126 102842
rect 35126 102790 35156 102842
rect 35180 102790 35190 102842
rect 35190 102790 35236 102842
rect 34940 102788 34996 102790
rect 35020 102788 35076 102790
rect 35100 102788 35156 102790
rect 35180 102788 35236 102790
rect 34940 101754 34996 101756
rect 35020 101754 35076 101756
rect 35100 101754 35156 101756
rect 35180 101754 35236 101756
rect 34940 101702 34986 101754
rect 34986 101702 34996 101754
rect 35020 101702 35050 101754
rect 35050 101702 35062 101754
rect 35062 101702 35076 101754
rect 35100 101702 35114 101754
rect 35114 101702 35126 101754
rect 35126 101702 35156 101754
rect 35180 101702 35190 101754
rect 35190 101702 35236 101754
rect 34940 101700 34996 101702
rect 35020 101700 35076 101702
rect 35100 101700 35156 101702
rect 35180 101700 35236 101702
rect 34940 100666 34996 100668
rect 35020 100666 35076 100668
rect 35100 100666 35156 100668
rect 35180 100666 35236 100668
rect 34940 100614 34986 100666
rect 34986 100614 34996 100666
rect 35020 100614 35050 100666
rect 35050 100614 35062 100666
rect 35062 100614 35076 100666
rect 35100 100614 35114 100666
rect 35114 100614 35126 100666
rect 35126 100614 35156 100666
rect 35180 100614 35190 100666
rect 35190 100614 35236 100666
rect 34940 100612 34996 100614
rect 35020 100612 35076 100614
rect 35100 100612 35156 100614
rect 35180 100612 35236 100614
rect 34940 99578 34996 99580
rect 35020 99578 35076 99580
rect 35100 99578 35156 99580
rect 35180 99578 35236 99580
rect 34940 99526 34986 99578
rect 34986 99526 34996 99578
rect 35020 99526 35050 99578
rect 35050 99526 35062 99578
rect 35062 99526 35076 99578
rect 35100 99526 35114 99578
rect 35114 99526 35126 99578
rect 35126 99526 35156 99578
rect 35180 99526 35190 99578
rect 35190 99526 35236 99578
rect 34940 99524 34996 99526
rect 35020 99524 35076 99526
rect 35100 99524 35156 99526
rect 35180 99524 35236 99526
rect 34940 98490 34996 98492
rect 35020 98490 35076 98492
rect 35100 98490 35156 98492
rect 35180 98490 35236 98492
rect 34940 98438 34986 98490
rect 34986 98438 34996 98490
rect 35020 98438 35050 98490
rect 35050 98438 35062 98490
rect 35062 98438 35076 98490
rect 35100 98438 35114 98490
rect 35114 98438 35126 98490
rect 35126 98438 35156 98490
rect 35180 98438 35190 98490
rect 35190 98438 35236 98490
rect 34940 98436 34996 98438
rect 35020 98436 35076 98438
rect 35100 98436 35156 98438
rect 35180 98436 35236 98438
rect 34940 97402 34996 97404
rect 35020 97402 35076 97404
rect 35100 97402 35156 97404
rect 35180 97402 35236 97404
rect 34940 97350 34986 97402
rect 34986 97350 34996 97402
rect 35020 97350 35050 97402
rect 35050 97350 35062 97402
rect 35062 97350 35076 97402
rect 35100 97350 35114 97402
rect 35114 97350 35126 97402
rect 35126 97350 35156 97402
rect 35180 97350 35190 97402
rect 35190 97350 35236 97402
rect 34940 97348 34996 97350
rect 35020 97348 35076 97350
rect 35100 97348 35156 97350
rect 35180 97348 35236 97350
rect 34940 96314 34996 96316
rect 35020 96314 35076 96316
rect 35100 96314 35156 96316
rect 35180 96314 35236 96316
rect 34940 96262 34986 96314
rect 34986 96262 34996 96314
rect 35020 96262 35050 96314
rect 35050 96262 35062 96314
rect 35062 96262 35076 96314
rect 35100 96262 35114 96314
rect 35114 96262 35126 96314
rect 35126 96262 35156 96314
rect 35180 96262 35190 96314
rect 35190 96262 35236 96314
rect 34940 96260 34996 96262
rect 35020 96260 35076 96262
rect 35100 96260 35156 96262
rect 35180 96260 35236 96262
rect 34940 95226 34996 95228
rect 35020 95226 35076 95228
rect 35100 95226 35156 95228
rect 35180 95226 35236 95228
rect 34940 95174 34986 95226
rect 34986 95174 34996 95226
rect 35020 95174 35050 95226
rect 35050 95174 35062 95226
rect 35062 95174 35076 95226
rect 35100 95174 35114 95226
rect 35114 95174 35126 95226
rect 35126 95174 35156 95226
rect 35180 95174 35190 95226
rect 35190 95174 35236 95226
rect 34940 95172 34996 95174
rect 35020 95172 35076 95174
rect 35100 95172 35156 95174
rect 35180 95172 35236 95174
rect 34940 94138 34996 94140
rect 35020 94138 35076 94140
rect 35100 94138 35156 94140
rect 35180 94138 35236 94140
rect 34940 94086 34986 94138
rect 34986 94086 34996 94138
rect 35020 94086 35050 94138
rect 35050 94086 35062 94138
rect 35062 94086 35076 94138
rect 35100 94086 35114 94138
rect 35114 94086 35126 94138
rect 35126 94086 35156 94138
rect 35180 94086 35190 94138
rect 35190 94086 35236 94138
rect 34940 94084 34996 94086
rect 35020 94084 35076 94086
rect 35100 94084 35156 94086
rect 35180 94084 35236 94086
rect 34940 93050 34996 93052
rect 35020 93050 35076 93052
rect 35100 93050 35156 93052
rect 35180 93050 35236 93052
rect 34940 92998 34986 93050
rect 34986 92998 34996 93050
rect 35020 92998 35050 93050
rect 35050 92998 35062 93050
rect 35062 92998 35076 93050
rect 35100 92998 35114 93050
rect 35114 92998 35126 93050
rect 35126 92998 35156 93050
rect 35180 92998 35190 93050
rect 35190 92998 35236 93050
rect 34940 92996 34996 92998
rect 35020 92996 35076 92998
rect 35100 92996 35156 92998
rect 35180 92996 35236 92998
rect 34940 91962 34996 91964
rect 35020 91962 35076 91964
rect 35100 91962 35156 91964
rect 35180 91962 35236 91964
rect 34940 91910 34986 91962
rect 34986 91910 34996 91962
rect 35020 91910 35050 91962
rect 35050 91910 35062 91962
rect 35062 91910 35076 91962
rect 35100 91910 35114 91962
rect 35114 91910 35126 91962
rect 35126 91910 35156 91962
rect 35180 91910 35190 91962
rect 35190 91910 35236 91962
rect 34940 91908 34996 91910
rect 35020 91908 35076 91910
rect 35100 91908 35156 91910
rect 35180 91908 35236 91910
rect 34940 90874 34996 90876
rect 35020 90874 35076 90876
rect 35100 90874 35156 90876
rect 35180 90874 35236 90876
rect 34940 90822 34986 90874
rect 34986 90822 34996 90874
rect 35020 90822 35050 90874
rect 35050 90822 35062 90874
rect 35062 90822 35076 90874
rect 35100 90822 35114 90874
rect 35114 90822 35126 90874
rect 35126 90822 35156 90874
rect 35180 90822 35190 90874
rect 35190 90822 35236 90874
rect 34940 90820 34996 90822
rect 35020 90820 35076 90822
rect 35100 90820 35156 90822
rect 35180 90820 35236 90822
rect 34940 89786 34996 89788
rect 35020 89786 35076 89788
rect 35100 89786 35156 89788
rect 35180 89786 35236 89788
rect 34940 89734 34986 89786
rect 34986 89734 34996 89786
rect 35020 89734 35050 89786
rect 35050 89734 35062 89786
rect 35062 89734 35076 89786
rect 35100 89734 35114 89786
rect 35114 89734 35126 89786
rect 35126 89734 35156 89786
rect 35180 89734 35190 89786
rect 35190 89734 35236 89786
rect 34940 89732 34996 89734
rect 35020 89732 35076 89734
rect 35100 89732 35156 89734
rect 35180 89732 35236 89734
rect 34940 88698 34996 88700
rect 35020 88698 35076 88700
rect 35100 88698 35156 88700
rect 35180 88698 35236 88700
rect 34940 88646 34986 88698
rect 34986 88646 34996 88698
rect 35020 88646 35050 88698
rect 35050 88646 35062 88698
rect 35062 88646 35076 88698
rect 35100 88646 35114 88698
rect 35114 88646 35126 88698
rect 35126 88646 35156 88698
rect 35180 88646 35190 88698
rect 35190 88646 35236 88698
rect 34940 88644 34996 88646
rect 35020 88644 35076 88646
rect 35100 88644 35156 88646
rect 35180 88644 35236 88646
rect 34940 87610 34996 87612
rect 35020 87610 35076 87612
rect 35100 87610 35156 87612
rect 35180 87610 35236 87612
rect 34940 87558 34986 87610
rect 34986 87558 34996 87610
rect 35020 87558 35050 87610
rect 35050 87558 35062 87610
rect 35062 87558 35076 87610
rect 35100 87558 35114 87610
rect 35114 87558 35126 87610
rect 35126 87558 35156 87610
rect 35180 87558 35190 87610
rect 35190 87558 35236 87610
rect 34940 87556 34996 87558
rect 35020 87556 35076 87558
rect 35100 87556 35156 87558
rect 35180 87556 35236 87558
rect 34940 86522 34996 86524
rect 35020 86522 35076 86524
rect 35100 86522 35156 86524
rect 35180 86522 35236 86524
rect 34940 86470 34986 86522
rect 34986 86470 34996 86522
rect 35020 86470 35050 86522
rect 35050 86470 35062 86522
rect 35062 86470 35076 86522
rect 35100 86470 35114 86522
rect 35114 86470 35126 86522
rect 35126 86470 35156 86522
rect 35180 86470 35190 86522
rect 35190 86470 35236 86522
rect 34940 86468 34996 86470
rect 35020 86468 35076 86470
rect 35100 86468 35156 86470
rect 35180 86468 35236 86470
rect 34940 85434 34996 85436
rect 35020 85434 35076 85436
rect 35100 85434 35156 85436
rect 35180 85434 35236 85436
rect 34940 85382 34986 85434
rect 34986 85382 34996 85434
rect 35020 85382 35050 85434
rect 35050 85382 35062 85434
rect 35062 85382 35076 85434
rect 35100 85382 35114 85434
rect 35114 85382 35126 85434
rect 35126 85382 35156 85434
rect 35180 85382 35190 85434
rect 35190 85382 35236 85434
rect 34940 85380 34996 85382
rect 35020 85380 35076 85382
rect 35100 85380 35156 85382
rect 35180 85380 35236 85382
rect 34940 84346 34996 84348
rect 35020 84346 35076 84348
rect 35100 84346 35156 84348
rect 35180 84346 35236 84348
rect 34940 84294 34986 84346
rect 34986 84294 34996 84346
rect 35020 84294 35050 84346
rect 35050 84294 35062 84346
rect 35062 84294 35076 84346
rect 35100 84294 35114 84346
rect 35114 84294 35126 84346
rect 35126 84294 35156 84346
rect 35180 84294 35190 84346
rect 35190 84294 35236 84346
rect 34940 84292 34996 84294
rect 35020 84292 35076 84294
rect 35100 84292 35156 84294
rect 35180 84292 35236 84294
rect 34940 83258 34996 83260
rect 35020 83258 35076 83260
rect 35100 83258 35156 83260
rect 35180 83258 35236 83260
rect 34940 83206 34986 83258
rect 34986 83206 34996 83258
rect 35020 83206 35050 83258
rect 35050 83206 35062 83258
rect 35062 83206 35076 83258
rect 35100 83206 35114 83258
rect 35114 83206 35126 83258
rect 35126 83206 35156 83258
rect 35180 83206 35190 83258
rect 35190 83206 35236 83258
rect 34940 83204 34996 83206
rect 35020 83204 35076 83206
rect 35100 83204 35156 83206
rect 35180 83204 35236 83206
rect 34940 82170 34996 82172
rect 35020 82170 35076 82172
rect 35100 82170 35156 82172
rect 35180 82170 35236 82172
rect 34940 82118 34986 82170
rect 34986 82118 34996 82170
rect 35020 82118 35050 82170
rect 35050 82118 35062 82170
rect 35062 82118 35076 82170
rect 35100 82118 35114 82170
rect 35114 82118 35126 82170
rect 35126 82118 35156 82170
rect 35180 82118 35190 82170
rect 35190 82118 35236 82170
rect 34940 82116 34996 82118
rect 35020 82116 35076 82118
rect 35100 82116 35156 82118
rect 35180 82116 35236 82118
rect 34940 81082 34996 81084
rect 35020 81082 35076 81084
rect 35100 81082 35156 81084
rect 35180 81082 35236 81084
rect 34940 81030 34986 81082
rect 34986 81030 34996 81082
rect 35020 81030 35050 81082
rect 35050 81030 35062 81082
rect 35062 81030 35076 81082
rect 35100 81030 35114 81082
rect 35114 81030 35126 81082
rect 35126 81030 35156 81082
rect 35180 81030 35190 81082
rect 35190 81030 35236 81082
rect 34940 81028 34996 81030
rect 35020 81028 35076 81030
rect 35100 81028 35156 81030
rect 35180 81028 35236 81030
rect 34940 79994 34996 79996
rect 35020 79994 35076 79996
rect 35100 79994 35156 79996
rect 35180 79994 35236 79996
rect 34940 79942 34986 79994
rect 34986 79942 34996 79994
rect 35020 79942 35050 79994
rect 35050 79942 35062 79994
rect 35062 79942 35076 79994
rect 35100 79942 35114 79994
rect 35114 79942 35126 79994
rect 35126 79942 35156 79994
rect 35180 79942 35190 79994
rect 35190 79942 35236 79994
rect 34940 79940 34996 79942
rect 35020 79940 35076 79942
rect 35100 79940 35156 79942
rect 35180 79940 35236 79942
rect 34940 78906 34996 78908
rect 35020 78906 35076 78908
rect 35100 78906 35156 78908
rect 35180 78906 35236 78908
rect 34940 78854 34986 78906
rect 34986 78854 34996 78906
rect 35020 78854 35050 78906
rect 35050 78854 35062 78906
rect 35062 78854 35076 78906
rect 35100 78854 35114 78906
rect 35114 78854 35126 78906
rect 35126 78854 35156 78906
rect 35180 78854 35190 78906
rect 35190 78854 35236 78906
rect 34940 78852 34996 78854
rect 35020 78852 35076 78854
rect 35100 78852 35156 78854
rect 35180 78852 35236 78854
rect 34940 77818 34996 77820
rect 35020 77818 35076 77820
rect 35100 77818 35156 77820
rect 35180 77818 35236 77820
rect 34940 77766 34986 77818
rect 34986 77766 34996 77818
rect 35020 77766 35050 77818
rect 35050 77766 35062 77818
rect 35062 77766 35076 77818
rect 35100 77766 35114 77818
rect 35114 77766 35126 77818
rect 35126 77766 35156 77818
rect 35180 77766 35190 77818
rect 35190 77766 35236 77818
rect 34940 77764 34996 77766
rect 35020 77764 35076 77766
rect 35100 77764 35156 77766
rect 35180 77764 35236 77766
rect 34940 76730 34996 76732
rect 35020 76730 35076 76732
rect 35100 76730 35156 76732
rect 35180 76730 35236 76732
rect 34940 76678 34986 76730
rect 34986 76678 34996 76730
rect 35020 76678 35050 76730
rect 35050 76678 35062 76730
rect 35062 76678 35076 76730
rect 35100 76678 35114 76730
rect 35114 76678 35126 76730
rect 35126 76678 35156 76730
rect 35180 76678 35190 76730
rect 35190 76678 35236 76730
rect 34940 76676 34996 76678
rect 35020 76676 35076 76678
rect 35100 76676 35156 76678
rect 35180 76676 35236 76678
rect 34940 75642 34996 75644
rect 35020 75642 35076 75644
rect 35100 75642 35156 75644
rect 35180 75642 35236 75644
rect 34940 75590 34986 75642
rect 34986 75590 34996 75642
rect 35020 75590 35050 75642
rect 35050 75590 35062 75642
rect 35062 75590 35076 75642
rect 35100 75590 35114 75642
rect 35114 75590 35126 75642
rect 35126 75590 35156 75642
rect 35180 75590 35190 75642
rect 35190 75590 35236 75642
rect 34940 75588 34996 75590
rect 35020 75588 35076 75590
rect 35100 75588 35156 75590
rect 35180 75588 35236 75590
rect 34940 74554 34996 74556
rect 35020 74554 35076 74556
rect 35100 74554 35156 74556
rect 35180 74554 35236 74556
rect 34940 74502 34986 74554
rect 34986 74502 34996 74554
rect 35020 74502 35050 74554
rect 35050 74502 35062 74554
rect 35062 74502 35076 74554
rect 35100 74502 35114 74554
rect 35114 74502 35126 74554
rect 35126 74502 35156 74554
rect 35180 74502 35190 74554
rect 35190 74502 35236 74554
rect 34940 74500 34996 74502
rect 35020 74500 35076 74502
rect 35100 74500 35156 74502
rect 35180 74500 35236 74502
rect 34940 73466 34996 73468
rect 35020 73466 35076 73468
rect 35100 73466 35156 73468
rect 35180 73466 35236 73468
rect 34940 73414 34986 73466
rect 34986 73414 34996 73466
rect 35020 73414 35050 73466
rect 35050 73414 35062 73466
rect 35062 73414 35076 73466
rect 35100 73414 35114 73466
rect 35114 73414 35126 73466
rect 35126 73414 35156 73466
rect 35180 73414 35190 73466
rect 35190 73414 35236 73466
rect 34940 73412 34996 73414
rect 35020 73412 35076 73414
rect 35100 73412 35156 73414
rect 35180 73412 35236 73414
rect 34940 72378 34996 72380
rect 35020 72378 35076 72380
rect 35100 72378 35156 72380
rect 35180 72378 35236 72380
rect 34940 72326 34986 72378
rect 34986 72326 34996 72378
rect 35020 72326 35050 72378
rect 35050 72326 35062 72378
rect 35062 72326 35076 72378
rect 35100 72326 35114 72378
rect 35114 72326 35126 72378
rect 35126 72326 35156 72378
rect 35180 72326 35190 72378
rect 35190 72326 35236 72378
rect 34940 72324 34996 72326
rect 35020 72324 35076 72326
rect 35100 72324 35156 72326
rect 35180 72324 35236 72326
rect 34940 71290 34996 71292
rect 35020 71290 35076 71292
rect 35100 71290 35156 71292
rect 35180 71290 35236 71292
rect 34940 71238 34986 71290
rect 34986 71238 34996 71290
rect 35020 71238 35050 71290
rect 35050 71238 35062 71290
rect 35062 71238 35076 71290
rect 35100 71238 35114 71290
rect 35114 71238 35126 71290
rect 35126 71238 35156 71290
rect 35180 71238 35190 71290
rect 35190 71238 35236 71290
rect 34940 71236 34996 71238
rect 35020 71236 35076 71238
rect 35100 71236 35156 71238
rect 35180 71236 35236 71238
rect 34940 70202 34996 70204
rect 35020 70202 35076 70204
rect 35100 70202 35156 70204
rect 35180 70202 35236 70204
rect 34940 70150 34986 70202
rect 34986 70150 34996 70202
rect 35020 70150 35050 70202
rect 35050 70150 35062 70202
rect 35062 70150 35076 70202
rect 35100 70150 35114 70202
rect 35114 70150 35126 70202
rect 35126 70150 35156 70202
rect 35180 70150 35190 70202
rect 35190 70150 35236 70202
rect 34940 70148 34996 70150
rect 35020 70148 35076 70150
rect 35100 70148 35156 70150
rect 35180 70148 35236 70150
rect 34940 69114 34996 69116
rect 35020 69114 35076 69116
rect 35100 69114 35156 69116
rect 35180 69114 35236 69116
rect 34940 69062 34986 69114
rect 34986 69062 34996 69114
rect 35020 69062 35050 69114
rect 35050 69062 35062 69114
rect 35062 69062 35076 69114
rect 35100 69062 35114 69114
rect 35114 69062 35126 69114
rect 35126 69062 35156 69114
rect 35180 69062 35190 69114
rect 35190 69062 35236 69114
rect 34940 69060 34996 69062
rect 35020 69060 35076 69062
rect 35100 69060 35156 69062
rect 35180 69060 35236 69062
rect 34940 68026 34996 68028
rect 35020 68026 35076 68028
rect 35100 68026 35156 68028
rect 35180 68026 35236 68028
rect 34940 67974 34986 68026
rect 34986 67974 34996 68026
rect 35020 67974 35050 68026
rect 35050 67974 35062 68026
rect 35062 67974 35076 68026
rect 35100 67974 35114 68026
rect 35114 67974 35126 68026
rect 35126 67974 35156 68026
rect 35180 67974 35190 68026
rect 35190 67974 35236 68026
rect 34940 67972 34996 67974
rect 35020 67972 35076 67974
rect 35100 67972 35156 67974
rect 35180 67972 35236 67974
rect 34940 66938 34996 66940
rect 35020 66938 35076 66940
rect 35100 66938 35156 66940
rect 35180 66938 35236 66940
rect 34940 66886 34986 66938
rect 34986 66886 34996 66938
rect 35020 66886 35050 66938
rect 35050 66886 35062 66938
rect 35062 66886 35076 66938
rect 35100 66886 35114 66938
rect 35114 66886 35126 66938
rect 35126 66886 35156 66938
rect 35180 66886 35190 66938
rect 35190 66886 35236 66938
rect 34940 66884 34996 66886
rect 35020 66884 35076 66886
rect 35100 66884 35156 66886
rect 35180 66884 35236 66886
rect 34940 65850 34996 65852
rect 35020 65850 35076 65852
rect 35100 65850 35156 65852
rect 35180 65850 35236 65852
rect 34940 65798 34986 65850
rect 34986 65798 34996 65850
rect 35020 65798 35050 65850
rect 35050 65798 35062 65850
rect 35062 65798 35076 65850
rect 35100 65798 35114 65850
rect 35114 65798 35126 65850
rect 35126 65798 35156 65850
rect 35180 65798 35190 65850
rect 35190 65798 35236 65850
rect 34940 65796 34996 65798
rect 35020 65796 35076 65798
rect 35100 65796 35156 65798
rect 35180 65796 35236 65798
rect 34940 64762 34996 64764
rect 35020 64762 35076 64764
rect 35100 64762 35156 64764
rect 35180 64762 35236 64764
rect 34940 64710 34986 64762
rect 34986 64710 34996 64762
rect 35020 64710 35050 64762
rect 35050 64710 35062 64762
rect 35062 64710 35076 64762
rect 35100 64710 35114 64762
rect 35114 64710 35126 64762
rect 35126 64710 35156 64762
rect 35180 64710 35190 64762
rect 35190 64710 35236 64762
rect 34940 64708 34996 64710
rect 35020 64708 35076 64710
rect 35100 64708 35156 64710
rect 35180 64708 35236 64710
rect 34940 63674 34996 63676
rect 35020 63674 35076 63676
rect 35100 63674 35156 63676
rect 35180 63674 35236 63676
rect 34940 63622 34986 63674
rect 34986 63622 34996 63674
rect 35020 63622 35050 63674
rect 35050 63622 35062 63674
rect 35062 63622 35076 63674
rect 35100 63622 35114 63674
rect 35114 63622 35126 63674
rect 35126 63622 35156 63674
rect 35180 63622 35190 63674
rect 35190 63622 35236 63674
rect 34940 63620 34996 63622
rect 35020 63620 35076 63622
rect 35100 63620 35156 63622
rect 35180 63620 35236 63622
rect 34940 62586 34996 62588
rect 35020 62586 35076 62588
rect 35100 62586 35156 62588
rect 35180 62586 35236 62588
rect 34940 62534 34986 62586
rect 34986 62534 34996 62586
rect 35020 62534 35050 62586
rect 35050 62534 35062 62586
rect 35062 62534 35076 62586
rect 35100 62534 35114 62586
rect 35114 62534 35126 62586
rect 35126 62534 35156 62586
rect 35180 62534 35190 62586
rect 35190 62534 35236 62586
rect 34940 62532 34996 62534
rect 35020 62532 35076 62534
rect 35100 62532 35156 62534
rect 35180 62532 35236 62534
rect 34940 61498 34996 61500
rect 35020 61498 35076 61500
rect 35100 61498 35156 61500
rect 35180 61498 35236 61500
rect 34940 61446 34986 61498
rect 34986 61446 34996 61498
rect 35020 61446 35050 61498
rect 35050 61446 35062 61498
rect 35062 61446 35076 61498
rect 35100 61446 35114 61498
rect 35114 61446 35126 61498
rect 35126 61446 35156 61498
rect 35180 61446 35190 61498
rect 35190 61446 35236 61498
rect 34940 61444 34996 61446
rect 35020 61444 35076 61446
rect 35100 61444 35156 61446
rect 35180 61444 35236 61446
rect 34940 60410 34996 60412
rect 35020 60410 35076 60412
rect 35100 60410 35156 60412
rect 35180 60410 35236 60412
rect 34940 60358 34986 60410
rect 34986 60358 34996 60410
rect 35020 60358 35050 60410
rect 35050 60358 35062 60410
rect 35062 60358 35076 60410
rect 35100 60358 35114 60410
rect 35114 60358 35126 60410
rect 35126 60358 35156 60410
rect 35180 60358 35190 60410
rect 35190 60358 35236 60410
rect 34940 60356 34996 60358
rect 35020 60356 35076 60358
rect 35100 60356 35156 60358
rect 35180 60356 35236 60358
rect 19580 59866 19636 59868
rect 19660 59866 19716 59868
rect 19740 59866 19796 59868
rect 19820 59866 19876 59868
rect 19580 59814 19626 59866
rect 19626 59814 19636 59866
rect 19660 59814 19690 59866
rect 19690 59814 19702 59866
rect 19702 59814 19716 59866
rect 19740 59814 19754 59866
rect 19754 59814 19766 59866
rect 19766 59814 19796 59866
rect 19820 59814 19830 59866
rect 19830 59814 19876 59866
rect 19580 59812 19636 59814
rect 19660 59812 19716 59814
rect 19740 59812 19796 59814
rect 19820 59812 19876 59814
rect 4220 59322 4276 59324
rect 4300 59322 4356 59324
rect 4380 59322 4436 59324
rect 4460 59322 4516 59324
rect 4220 59270 4266 59322
rect 4266 59270 4276 59322
rect 4300 59270 4330 59322
rect 4330 59270 4342 59322
rect 4342 59270 4356 59322
rect 4380 59270 4394 59322
rect 4394 59270 4406 59322
rect 4406 59270 4436 59322
rect 4460 59270 4470 59322
rect 4470 59270 4516 59322
rect 4220 59268 4276 59270
rect 4300 59268 4356 59270
rect 4380 59268 4436 59270
rect 4460 59268 4516 59270
rect 4220 58234 4276 58236
rect 4300 58234 4356 58236
rect 4380 58234 4436 58236
rect 4460 58234 4516 58236
rect 4220 58182 4266 58234
rect 4266 58182 4276 58234
rect 4300 58182 4330 58234
rect 4330 58182 4342 58234
rect 4342 58182 4356 58234
rect 4380 58182 4394 58234
rect 4394 58182 4406 58234
rect 4406 58182 4436 58234
rect 4460 58182 4470 58234
rect 4470 58182 4516 58234
rect 4220 58180 4276 58182
rect 4300 58180 4356 58182
rect 4380 58180 4436 58182
rect 4460 58180 4516 58182
rect 4220 57146 4276 57148
rect 4300 57146 4356 57148
rect 4380 57146 4436 57148
rect 4460 57146 4516 57148
rect 4220 57094 4266 57146
rect 4266 57094 4276 57146
rect 4300 57094 4330 57146
rect 4330 57094 4342 57146
rect 4342 57094 4356 57146
rect 4380 57094 4394 57146
rect 4394 57094 4406 57146
rect 4406 57094 4436 57146
rect 4460 57094 4470 57146
rect 4470 57094 4516 57146
rect 4220 57092 4276 57094
rect 4300 57092 4356 57094
rect 4380 57092 4436 57094
rect 4460 57092 4516 57094
rect 4220 56058 4276 56060
rect 4300 56058 4356 56060
rect 4380 56058 4436 56060
rect 4460 56058 4516 56060
rect 4220 56006 4266 56058
rect 4266 56006 4276 56058
rect 4300 56006 4330 56058
rect 4330 56006 4342 56058
rect 4342 56006 4356 56058
rect 4380 56006 4394 56058
rect 4394 56006 4406 56058
rect 4406 56006 4436 56058
rect 4460 56006 4470 56058
rect 4470 56006 4516 56058
rect 4220 56004 4276 56006
rect 4300 56004 4356 56006
rect 4380 56004 4436 56006
rect 4460 56004 4516 56006
rect 4220 54970 4276 54972
rect 4300 54970 4356 54972
rect 4380 54970 4436 54972
rect 4460 54970 4516 54972
rect 4220 54918 4266 54970
rect 4266 54918 4276 54970
rect 4300 54918 4330 54970
rect 4330 54918 4342 54970
rect 4342 54918 4356 54970
rect 4380 54918 4394 54970
rect 4394 54918 4406 54970
rect 4406 54918 4436 54970
rect 4460 54918 4470 54970
rect 4470 54918 4516 54970
rect 4220 54916 4276 54918
rect 4300 54916 4356 54918
rect 4380 54916 4436 54918
rect 4460 54916 4516 54918
rect 4220 53882 4276 53884
rect 4300 53882 4356 53884
rect 4380 53882 4436 53884
rect 4460 53882 4516 53884
rect 4220 53830 4266 53882
rect 4266 53830 4276 53882
rect 4300 53830 4330 53882
rect 4330 53830 4342 53882
rect 4342 53830 4356 53882
rect 4380 53830 4394 53882
rect 4394 53830 4406 53882
rect 4406 53830 4436 53882
rect 4460 53830 4470 53882
rect 4470 53830 4516 53882
rect 4220 53828 4276 53830
rect 4300 53828 4356 53830
rect 4380 53828 4436 53830
rect 4460 53828 4516 53830
rect 4220 52794 4276 52796
rect 4300 52794 4356 52796
rect 4380 52794 4436 52796
rect 4460 52794 4516 52796
rect 4220 52742 4266 52794
rect 4266 52742 4276 52794
rect 4300 52742 4330 52794
rect 4330 52742 4342 52794
rect 4342 52742 4356 52794
rect 4380 52742 4394 52794
rect 4394 52742 4406 52794
rect 4406 52742 4436 52794
rect 4460 52742 4470 52794
rect 4470 52742 4516 52794
rect 4220 52740 4276 52742
rect 4300 52740 4356 52742
rect 4380 52740 4436 52742
rect 4460 52740 4516 52742
rect 4220 51706 4276 51708
rect 4300 51706 4356 51708
rect 4380 51706 4436 51708
rect 4460 51706 4516 51708
rect 4220 51654 4266 51706
rect 4266 51654 4276 51706
rect 4300 51654 4330 51706
rect 4330 51654 4342 51706
rect 4342 51654 4356 51706
rect 4380 51654 4394 51706
rect 4394 51654 4406 51706
rect 4406 51654 4436 51706
rect 4460 51654 4470 51706
rect 4470 51654 4516 51706
rect 4220 51652 4276 51654
rect 4300 51652 4356 51654
rect 4380 51652 4436 51654
rect 4460 51652 4516 51654
rect 4220 50618 4276 50620
rect 4300 50618 4356 50620
rect 4380 50618 4436 50620
rect 4460 50618 4516 50620
rect 4220 50566 4266 50618
rect 4266 50566 4276 50618
rect 4300 50566 4330 50618
rect 4330 50566 4342 50618
rect 4342 50566 4356 50618
rect 4380 50566 4394 50618
rect 4394 50566 4406 50618
rect 4406 50566 4436 50618
rect 4460 50566 4470 50618
rect 4470 50566 4516 50618
rect 4220 50564 4276 50566
rect 4300 50564 4356 50566
rect 4380 50564 4436 50566
rect 4460 50564 4516 50566
rect 4220 49530 4276 49532
rect 4300 49530 4356 49532
rect 4380 49530 4436 49532
rect 4460 49530 4516 49532
rect 4220 49478 4266 49530
rect 4266 49478 4276 49530
rect 4300 49478 4330 49530
rect 4330 49478 4342 49530
rect 4342 49478 4356 49530
rect 4380 49478 4394 49530
rect 4394 49478 4406 49530
rect 4406 49478 4436 49530
rect 4460 49478 4470 49530
rect 4470 49478 4516 49530
rect 4220 49476 4276 49478
rect 4300 49476 4356 49478
rect 4380 49476 4436 49478
rect 4460 49476 4516 49478
rect 4220 48442 4276 48444
rect 4300 48442 4356 48444
rect 4380 48442 4436 48444
rect 4460 48442 4516 48444
rect 4220 48390 4266 48442
rect 4266 48390 4276 48442
rect 4300 48390 4330 48442
rect 4330 48390 4342 48442
rect 4342 48390 4356 48442
rect 4380 48390 4394 48442
rect 4394 48390 4406 48442
rect 4406 48390 4436 48442
rect 4460 48390 4470 48442
rect 4470 48390 4516 48442
rect 4220 48388 4276 48390
rect 4300 48388 4356 48390
rect 4380 48388 4436 48390
rect 4460 48388 4516 48390
rect 4220 47354 4276 47356
rect 4300 47354 4356 47356
rect 4380 47354 4436 47356
rect 4460 47354 4516 47356
rect 4220 47302 4266 47354
rect 4266 47302 4276 47354
rect 4300 47302 4330 47354
rect 4330 47302 4342 47354
rect 4342 47302 4356 47354
rect 4380 47302 4394 47354
rect 4394 47302 4406 47354
rect 4406 47302 4436 47354
rect 4460 47302 4470 47354
rect 4470 47302 4516 47354
rect 4220 47300 4276 47302
rect 4300 47300 4356 47302
rect 4380 47300 4436 47302
rect 4460 47300 4516 47302
rect 4220 46266 4276 46268
rect 4300 46266 4356 46268
rect 4380 46266 4436 46268
rect 4460 46266 4516 46268
rect 4220 46214 4266 46266
rect 4266 46214 4276 46266
rect 4300 46214 4330 46266
rect 4330 46214 4342 46266
rect 4342 46214 4356 46266
rect 4380 46214 4394 46266
rect 4394 46214 4406 46266
rect 4406 46214 4436 46266
rect 4460 46214 4470 46266
rect 4470 46214 4516 46266
rect 4220 46212 4276 46214
rect 4300 46212 4356 46214
rect 4380 46212 4436 46214
rect 4460 46212 4516 46214
rect 4220 45178 4276 45180
rect 4300 45178 4356 45180
rect 4380 45178 4436 45180
rect 4460 45178 4516 45180
rect 4220 45126 4266 45178
rect 4266 45126 4276 45178
rect 4300 45126 4330 45178
rect 4330 45126 4342 45178
rect 4342 45126 4356 45178
rect 4380 45126 4394 45178
rect 4394 45126 4406 45178
rect 4406 45126 4436 45178
rect 4460 45126 4470 45178
rect 4470 45126 4516 45178
rect 4220 45124 4276 45126
rect 4300 45124 4356 45126
rect 4380 45124 4436 45126
rect 4460 45124 4516 45126
rect 4220 44090 4276 44092
rect 4300 44090 4356 44092
rect 4380 44090 4436 44092
rect 4460 44090 4516 44092
rect 4220 44038 4266 44090
rect 4266 44038 4276 44090
rect 4300 44038 4330 44090
rect 4330 44038 4342 44090
rect 4342 44038 4356 44090
rect 4380 44038 4394 44090
rect 4394 44038 4406 44090
rect 4406 44038 4436 44090
rect 4460 44038 4470 44090
rect 4470 44038 4516 44090
rect 4220 44036 4276 44038
rect 4300 44036 4356 44038
rect 4380 44036 4436 44038
rect 4460 44036 4516 44038
rect 4220 43002 4276 43004
rect 4300 43002 4356 43004
rect 4380 43002 4436 43004
rect 4460 43002 4516 43004
rect 4220 42950 4266 43002
rect 4266 42950 4276 43002
rect 4300 42950 4330 43002
rect 4330 42950 4342 43002
rect 4342 42950 4356 43002
rect 4380 42950 4394 43002
rect 4394 42950 4406 43002
rect 4406 42950 4436 43002
rect 4460 42950 4470 43002
rect 4470 42950 4516 43002
rect 4220 42948 4276 42950
rect 4300 42948 4356 42950
rect 4380 42948 4436 42950
rect 4460 42948 4516 42950
rect 4220 41914 4276 41916
rect 4300 41914 4356 41916
rect 4380 41914 4436 41916
rect 4460 41914 4516 41916
rect 4220 41862 4266 41914
rect 4266 41862 4276 41914
rect 4300 41862 4330 41914
rect 4330 41862 4342 41914
rect 4342 41862 4356 41914
rect 4380 41862 4394 41914
rect 4394 41862 4406 41914
rect 4406 41862 4436 41914
rect 4460 41862 4470 41914
rect 4470 41862 4516 41914
rect 4220 41860 4276 41862
rect 4300 41860 4356 41862
rect 4380 41860 4436 41862
rect 4460 41860 4516 41862
rect 4220 40826 4276 40828
rect 4300 40826 4356 40828
rect 4380 40826 4436 40828
rect 4460 40826 4516 40828
rect 4220 40774 4266 40826
rect 4266 40774 4276 40826
rect 4300 40774 4330 40826
rect 4330 40774 4342 40826
rect 4342 40774 4356 40826
rect 4380 40774 4394 40826
rect 4394 40774 4406 40826
rect 4406 40774 4436 40826
rect 4460 40774 4470 40826
rect 4470 40774 4516 40826
rect 4220 40772 4276 40774
rect 4300 40772 4356 40774
rect 4380 40772 4436 40774
rect 4460 40772 4516 40774
rect 4220 39738 4276 39740
rect 4300 39738 4356 39740
rect 4380 39738 4436 39740
rect 4460 39738 4516 39740
rect 4220 39686 4266 39738
rect 4266 39686 4276 39738
rect 4300 39686 4330 39738
rect 4330 39686 4342 39738
rect 4342 39686 4356 39738
rect 4380 39686 4394 39738
rect 4394 39686 4406 39738
rect 4406 39686 4436 39738
rect 4460 39686 4470 39738
rect 4470 39686 4516 39738
rect 4220 39684 4276 39686
rect 4300 39684 4356 39686
rect 4380 39684 4436 39686
rect 4460 39684 4516 39686
rect 4220 38650 4276 38652
rect 4300 38650 4356 38652
rect 4380 38650 4436 38652
rect 4460 38650 4516 38652
rect 4220 38598 4266 38650
rect 4266 38598 4276 38650
rect 4300 38598 4330 38650
rect 4330 38598 4342 38650
rect 4342 38598 4356 38650
rect 4380 38598 4394 38650
rect 4394 38598 4406 38650
rect 4406 38598 4436 38650
rect 4460 38598 4470 38650
rect 4470 38598 4516 38650
rect 4220 38596 4276 38598
rect 4300 38596 4356 38598
rect 4380 38596 4436 38598
rect 4460 38596 4516 38598
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 19580 58778 19636 58780
rect 19660 58778 19716 58780
rect 19740 58778 19796 58780
rect 19820 58778 19876 58780
rect 19580 58726 19626 58778
rect 19626 58726 19636 58778
rect 19660 58726 19690 58778
rect 19690 58726 19702 58778
rect 19702 58726 19716 58778
rect 19740 58726 19754 58778
rect 19754 58726 19766 58778
rect 19766 58726 19796 58778
rect 19820 58726 19830 58778
rect 19830 58726 19876 58778
rect 19580 58724 19636 58726
rect 19660 58724 19716 58726
rect 19740 58724 19796 58726
rect 19820 58724 19876 58726
rect 19580 57690 19636 57692
rect 19660 57690 19716 57692
rect 19740 57690 19796 57692
rect 19820 57690 19876 57692
rect 19580 57638 19626 57690
rect 19626 57638 19636 57690
rect 19660 57638 19690 57690
rect 19690 57638 19702 57690
rect 19702 57638 19716 57690
rect 19740 57638 19754 57690
rect 19754 57638 19766 57690
rect 19766 57638 19796 57690
rect 19820 57638 19830 57690
rect 19830 57638 19876 57690
rect 19580 57636 19636 57638
rect 19660 57636 19716 57638
rect 19740 57636 19796 57638
rect 19820 57636 19876 57638
rect 19580 56602 19636 56604
rect 19660 56602 19716 56604
rect 19740 56602 19796 56604
rect 19820 56602 19876 56604
rect 19580 56550 19626 56602
rect 19626 56550 19636 56602
rect 19660 56550 19690 56602
rect 19690 56550 19702 56602
rect 19702 56550 19716 56602
rect 19740 56550 19754 56602
rect 19754 56550 19766 56602
rect 19766 56550 19796 56602
rect 19820 56550 19830 56602
rect 19830 56550 19876 56602
rect 19580 56548 19636 56550
rect 19660 56548 19716 56550
rect 19740 56548 19796 56550
rect 19820 56548 19876 56550
rect 19580 55514 19636 55516
rect 19660 55514 19716 55516
rect 19740 55514 19796 55516
rect 19820 55514 19876 55516
rect 19580 55462 19626 55514
rect 19626 55462 19636 55514
rect 19660 55462 19690 55514
rect 19690 55462 19702 55514
rect 19702 55462 19716 55514
rect 19740 55462 19754 55514
rect 19754 55462 19766 55514
rect 19766 55462 19796 55514
rect 19820 55462 19830 55514
rect 19830 55462 19876 55514
rect 19580 55460 19636 55462
rect 19660 55460 19716 55462
rect 19740 55460 19796 55462
rect 19820 55460 19876 55462
rect 19580 54426 19636 54428
rect 19660 54426 19716 54428
rect 19740 54426 19796 54428
rect 19820 54426 19876 54428
rect 19580 54374 19626 54426
rect 19626 54374 19636 54426
rect 19660 54374 19690 54426
rect 19690 54374 19702 54426
rect 19702 54374 19716 54426
rect 19740 54374 19754 54426
rect 19754 54374 19766 54426
rect 19766 54374 19796 54426
rect 19820 54374 19830 54426
rect 19830 54374 19876 54426
rect 19580 54372 19636 54374
rect 19660 54372 19716 54374
rect 19740 54372 19796 54374
rect 19820 54372 19876 54374
rect 19580 53338 19636 53340
rect 19660 53338 19716 53340
rect 19740 53338 19796 53340
rect 19820 53338 19876 53340
rect 19580 53286 19626 53338
rect 19626 53286 19636 53338
rect 19660 53286 19690 53338
rect 19690 53286 19702 53338
rect 19702 53286 19716 53338
rect 19740 53286 19754 53338
rect 19754 53286 19766 53338
rect 19766 53286 19796 53338
rect 19820 53286 19830 53338
rect 19830 53286 19876 53338
rect 19580 53284 19636 53286
rect 19660 53284 19716 53286
rect 19740 53284 19796 53286
rect 19820 53284 19876 53286
rect 19580 52250 19636 52252
rect 19660 52250 19716 52252
rect 19740 52250 19796 52252
rect 19820 52250 19876 52252
rect 19580 52198 19626 52250
rect 19626 52198 19636 52250
rect 19660 52198 19690 52250
rect 19690 52198 19702 52250
rect 19702 52198 19716 52250
rect 19740 52198 19754 52250
rect 19754 52198 19766 52250
rect 19766 52198 19796 52250
rect 19820 52198 19830 52250
rect 19830 52198 19876 52250
rect 19580 52196 19636 52198
rect 19660 52196 19716 52198
rect 19740 52196 19796 52198
rect 19820 52196 19876 52198
rect 19580 51162 19636 51164
rect 19660 51162 19716 51164
rect 19740 51162 19796 51164
rect 19820 51162 19876 51164
rect 19580 51110 19626 51162
rect 19626 51110 19636 51162
rect 19660 51110 19690 51162
rect 19690 51110 19702 51162
rect 19702 51110 19716 51162
rect 19740 51110 19754 51162
rect 19754 51110 19766 51162
rect 19766 51110 19796 51162
rect 19820 51110 19830 51162
rect 19830 51110 19876 51162
rect 19580 51108 19636 51110
rect 19660 51108 19716 51110
rect 19740 51108 19796 51110
rect 19820 51108 19876 51110
rect 19580 50074 19636 50076
rect 19660 50074 19716 50076
rect 19740 50074 19796 50076
rect 19820 50074 19876 50076
rect 19580 50022 19626 50074
rect 19626 50022 19636 50074
rect 19660 50022 19690 50074
rect 19690 50022 19702 50074
rect 19702 50022 19716 50074
rect 19740 50022 19754 50074
rect 19754 50022 19766 50074
rect 19766 50022 19796 50074
rect 19820 50022 19830 50074
rect 19830 50022 19876 50074
rect 19580 50020 19636 50022
rect 19660 50020 19716 50022
rect 19740 50020 19796 50022
rect 19820 50020 19876 50022
rect 19580 48986 19636 48988
rect 19660 48986 19716 48988
rect 19740 48986 19796 48988
rect 19820 48986 19876 48988
rect 19580 48934 19626 48986
rect 19626 48934 19636 48986
rect 19660 48934 19690 48986
rect 19690 48934 19702 48986
rect 19702 48934 19716 48986
rect 19740 48934 19754 48986
rect 19754 48934 19766 48986
rect 19766 48934 19796 48986
rect 19820 48934 19830 48986
rect 19830 48934 19876 48986
rect 19580 48932 19636 48934
rect 19660 48932 19716 48934
rect 19740 48932 19796 48934
rect 19820 48932 19876 48934
rect 19580 47898 19636 47900
rect 19660 47898 19716 47900
rect 19740 47898 19796 47900
rect 19820 47898 19876 47900
rect 19580 47846 19626 47898
rect 19626 47846 19636 47898
rect 19660 47846 19690 47898
rect 19690 47846 19702 47898
rect 19702 47846 19716 47898
rect 19740 47846 19754 47898
rect 19754 47846 19766 47898
rect 19766 47846 19796 47898
rect 19820 47846 19830 47898
rect 19830 47846 19876 47898
rect 19580 47844 19636 47846
rect 19660 47844 19716 47846
rect 19740 47844 19796 47846
rect 19820 47844 19876 47846
rect 19580 46810 19636 46812
rect 19660 46810 19716 46812
rect 19740 46810 19796 46812
rect 19820 46810 19876 46812
rect 19580 46758 19626 46810
rect 19626 46758 19636 46810
rect 19660 46758 19690 46810
rect 19690 46758 19702 46810
rect 19702 46758 19716 46810
rect 19740 46758 19754 46810
rect 19754 46758 19766 46810
rect 19766 46758 19796 46810
rect 19820 46758 19830 46810
rect 19830 46758 19876 46810
rect 19580 46756 19636 46758
rect 19660 46756 19716 46758
rect 19740 46756 19796 46758
rect 19820 46756 19876 46758
rect 19580 45722 19636 45724
rect 19660 45722 19716 45724
rect 19740 45722 19796 45724
rect 19820 45722 19876 45724
rect 19580 45670 19626 45722
rect 19626 45670 19636 45722
rect 19660 45670 19690 45722
rect 19690 45670 19702 45722
rect 19702 45670 19716 45722
rect 19740 45670 19754 45722
rect 19754 45670 19766 45722
rect 19766 45670 19796 45722
rect 19820 45670 19830 45722
rect 19830 45670 19876 45722
rect 19580 45668 19636 45670
rect 19660 45668 19716 45670
rect 19740 45668 19796 45670
rect 19820 45668 19876 45670
rect 19580 44634 19636 44636
rect 19660 44634 19716 44636
rect 19740 44634 19796 44636
rect 19820 44634 19876 44636
rect 19580 44582 19626 44634
rect 19626 44582 19636 44634
rect 19660 44582 19690 44634
rect 19690 44582 19702 44634
rect 19702 44582 19716 44634
rect 19740 44582 19754 44634
rect 19754 44582 19766 44634
rect 19766 44582 19796 44634
rect 19820 44582 19830 44634
rect 19830 44582 19876 44634
rect 19580 44580 19636 44582
rect 19660 44580 19716 44582
rect 19740 44580 19796 44582
rect 19820 44580 19876 44582
rect 19580 43546 19636 43548
rect 19660 43546 19716 43548
rect 19740 43546 19796 43548
rect 19820 43546 19876 43548
rect 19580 43494 19626 43546
rect 19626 43494 19636 43546
rect 19660 43494 19690 43546
rect 19690 43494 19702 43546
rect 19702 43494 19716 43546
rect 19740 43494 19754 43546
rect 19754 43494 19766 43546
rect 19766 43494 19796 43546
rect 19820 43494 19830 43546
rect 19830 43494 19876 43546
rect 19580 43492 19636 43494
rect 19660 43492 19716 43494
rect 19740 43492 19796 43494
rect 19820 43492 19876 43494
rect 19580 42458 19636 42460
rect 19660 42458 19716 42460
rect 19740 42458 19796 42460
rect 19820 42458 19876 42460
rect 19580 42406 19626 42458
rect 19626 42406 19636 42458
rect 19660 42406 19690 42458
rect 19690 42406 19702 42458
rect 19702 42406 19716 42458
rect 19740 42406 19754 42458
rect 19754 42406 19766 42458
rect 19766 42406 19796 42458
rect 19820 42406 19830 42458
rect 19830 42406 19876 42458
rect 19580 42404 19636 42406
rect 19660 42404 19716 42406
rect 19740 42404 19796 42406
rect 19820 42404 19876 42406
rect 19580 41370 19636 41372
rect 19660 41370 19716 41372
rect 19740 41370 19796 41372
rect 19820 41370 19876 41372
rect 19580 41318 19626 41370
rect 19626 41318 19636 41370
rect 19660 41318 19690 41370
rect 19690 41318 19702 41370
rect 19702 41318 19716 41370
rect 19740 41318 19754 41370
rect 19754 41318 19766 41370
rect 19766 41318 19796 41370
rect 19820 41318 19830 41370
rect 19830 41318 19876 41370
rect 19580 41316 19636 41318
rect 19660 41316 19716 41318
rect 19740 41316 19796 41318
rect 19820 41316 19876 41318
rect 19580 40282 19636 40284
rect 19660 40282 19716 40284
rect 19740 40282 19796 40284
rect 19820 40282 19876 40284
rect 19580 40230 19626 40282
rect 19626 40230 19636 40282
rect 19660 40230 19690 40282
rect 19690 40230 19702 40282
rect 19702 40230 19716 40282
rect 19740 40230 19754 40282
rect 19754 40230 19766 40282
rect 19766 40230 19796 40282
rect 19820 40230 19830 40282
rect 19830 40230 19876 40282
rect 19580 40228 19636 40230
rect 19660 40228 19716 40230
rect 19740 40228 19796 40230
rect 19820 40228 19876 40230
rect 19580 39194 19636 39196
rect 19660 39194 19716 39196
rect 19740 39194 19796 39196
rect 19820 39194 19876 39196
rect 19580 39142 19626 39194
rect 19626 39142 19636 39194
rect 19660 39142 19690 39194
rect 19690 39142 19702 39194
rect 19702 39142 19716 39194
rect 19740 39142 19754 39194
rect 19754 39142 19766 39194
rect 19766 39142 19796 39194
rect 19820 39142 19830 39194
rect 19830 39142 19876 39194
rect 19580 39140 19636 39142
rect 19660 39140 19716 39142
rect 19740 39140 19796 39142
rect 19820 39140 19876 39142
rect 19580 38106 19636 38108
rect 19660 38106 19716 38108
rect 19740 38106 19796 38108
rect 19820 38106 19876 38108
rect 19580 38054 19626 38106
rect 19626 38054 19636 38106
rect 19660 38054 19690 38106
rect 19690 38054 19702 38106
rect 19702 38054 19716 38106
rect 19740 38054 19754 38106
rect 19754 38054 19766 38106
rect 19766 38054 19796 38106
rect 19820 38054 19830 38106
rect 19830 38054 19876 38106
rect 19580 38052 19636 38054
rect 19660 38052 19716 38054
rect 19740 38052 19796 38054
rect 19820 38052 19876 38054
rect 19580 37018 19636 37020
rect 19660 37018 19716 37020
rect 19740 37018 19796 37020
rect 19820 37018 19876 37020
rect 19580 36966 19626 37018
rect 19626 36966 19636 37018
rect 19660 36966 19690 37018
rect 19690 36966 19702 37018
rect 19702 36966 19716 37018
rect 19740 36966 19754 37018
rect 19754 36966 19766 37018
rect 19766 36966 19796 37018
rect 19820 36966 19830 37018
rect 19830 36966 19876 37018
rect 19580 36964 19636 36966
rect 19660 36964 19716 36966
rect 19740 36964 19796 36966
rect 19820 36964 19876 36966
rect 19580 35930 19636 35932
rect 19660 35930 19716 35932
rect 19740 35930 19796 35932
rect 19820 35930 19876 35932
rect 19580 35878 19626 35930
rect 19626 35878 19636 35930
rect 19660 35878 19690 35930
rect 19690 35878 19702 35930
rect 19702 35878 19716 35930
rect 19740 35878 19754 35930
rect 19754 35878 19766 35930
rect 19766 35878 19796 35930
rect 19820 35878 19830 35930
rect 19830 35878 19876 35930
rect 19580 35876 19636 35878
rect 19660 35876 19716 35878
rect 19740 35876 19796 35878
rect 19820 35876 19876 35878
rect 19580 34842 19636 34844
rect 19660 34842 19716 34844
rect 19740 34842 19796 34844
rect 19820 34842 19876 34844
rect 19580 34790 19626 34842
rect 19626 34790 19636 34842
rect 19660 34790 19690 34842
rect 19690 34790 19702 34842
rect 19702 34790 19716 34842
rect 19740 34790 19754 34842
rect 19754 34790 19766 34842
rect 19766 34790 19796 34842
rect 19820 34790 19830 34842
rect 19830 34790 19876 34842
rect 19580 34788 19636 34790
rect 19660 34788 19716 34790
rect 19740 34788 19796 34790
rect 19820 34788 19876 34790
rect 19580 33754 19636 33756
rect 19660 33754 19716 33756
rect 19740 33754 19796 33756
rect 19820 33754 19876 33756
rect 19580 33702 19626 33754
rect 19626 33702 19636 33754
rect 19660 33702 19690 33754
rect 19690 33702 19702 33754
rect 19702 33702 19716 33754
rect 19740 33702 19754 33754
rect 19754 33702 19766 33754
rect 19766 33702 19796 33754
rect 19820 33702 19830 33754
rect 19830 33702 19876 33754
rect 19580 33700 19636 33702
rect 19660 33700 19716 33702
rect 19740 33700 19796 33702
rect 19820 33700 19876 33702
rect 19580 32666 19636 32668
rect 19660 32666 19716 32668
rect 19740 32666 19796 32668
rect 19820 32666 19876 32668
rect 19580 32614 19626 32666
rect 19626 32614 19636 32666
rect 19660 32614 19690 32666
rect 19690 32614 19702 32666
rect 19702 32614 19716 32666
rect 19740 32614 19754 32666
rect 19754 32614 19766 32666
rect 19766 32614 19796 32666
rect 19820 32614 19830 32666
rect 19830 32614 19876 32666
rect 19580 32612 19636 32614
rect 19660 32612 19716 32614
rect 19740 32612 19796 32614
rect 19820 32612 19876 32614
rect 19580 31578 19636 31580
rect 19660 31578 19716 31580
rect 19740 31578 19796 31580
rect 19820 31578 19876 31580
rect 19580 31526 19626 31578
rect 19626 31526 19636 31578
rect 19660 31526 19690 31578
rect 19690 31526 19702 31578
rect 19702 31526 19716 31578
rect 19740 31526 19754 31578
rect 19754 31526 19766 31578
rect 19766 31526 19796 31578
rect 19820 31526 19830 31578
rect 19830 31526 19876 31578
rect 19580 31524 19636 31526
rect 19660 31524 19716 31526
rect 19740 31524 19796 31526
rect 19820 31524 19876 31526
rect 19580 30490 19636 30492
rect 19660 30490 19716 30492
rect 19740 30490 19796 30492
rect 19820 30490 19876 30492
rect 19580 30438 19626 30490
rect 19626 30438 19636 30490
rect 19660 30438 19690 30490
rect 19690 30438 19702 30490
rect 19702 30438 19716 30490
rect 19740 30438 19754 30490
rect 19754 30438 19766 30490
rect 19766 30438 19796 30490
rect 19820 30438 19830 30490
rect 19830 30438 19876 30490
rect 19580 30436 19636 30438
rect 19660 30436 19716 30438
rect 19740 30436 19796 30438
rect 19820 30436 19876 30438
rect 19580 29402 19636 29404
rect 19660 29402 19716 29404
rect 19740 29402 19796 29404
rect 19820 29402 19876 29404
rect 19580 29350 19626 29402
rect 19626 29350 19636 29402
rect 19660 29350 19690 29402
rect 19690 29350 19702 29402
rect 19702 29350 19716 29402
rect 19740 29350 19754 29402
rect 19754 29350 19766 29402
rect 19766 29350 19796 29402
rect 19820 29350 19830 29402
rect 19830 29350 19876 29402
rect 19580 29348 19636 29350
rect 19660 29348 19716 29350
rect 19740 29348 19796 29350
rect 19820 29348 19876 29350
rect 19580 28314 19636 28316
rect 19660 28314 19716 28316
rect 19740 28314 19796 28316
rect 19820 28314 19876 28316
rect 19580 28262 19626 28314
rect 19626 28262 19636 28314
rect 19660 28262 19690 28314
rect 19690 28262 19702 28314
rect 19702 28262 19716 28314
rect 19740 28262 19754 28314
rect 19754 28262 19766 28314
rect 19766 28262 19796 28314
rect 19820 28262 19830 28314
rect 19830 28262 19876 28314
rect 19580 28260 19636 28262
rect 19660 28260 19716 28262
rect 19740 28260 19796 28262
rect 19820 28260 19876 28262
rect 19580 27226 19636 27228
rect 19660 27226 19716 27228
rect 19740 27226 19796 27228
rect 19820 27226 19876 27228
rect 19580 27174 19626 27226
rect 19626 27174 19636 27226
rect 19660 27174 19690 27226
rect 19690 27174 19702 27226
rect 19702 27174 19716 27226
rect 19740 27174 19754 27226
rect 19754 27174 19766 27226
rect 19766 27174 19796 27226
rect 19820 27174 19830 27226
rect 19830 27174 19876 27226
rect 19580 27172 19636 27174
rect 19660 27172 19716 27174
rect 19740 27172 19796 27174
rect 19820 27172 19876 27174
rect 19580 26138 19636 26140
rect 19660 26138 19716 26140
rect 19740 26138 19796 26140
rect 19820 26138 19876 26140
rect 19580 26086 19626 26138
rect 19626 26086 19636 26138
rect 19660 26086 19690 26138
rect 19690 26086 19702 26138
rect 19702 26086 19716 26138
rect 19740 26086 19754 26138
rect 19754 26086 19766 26138
rect 19766 26086 19796 26138
rect 19820 26086 19830 26138
rect 19830 26086 19876 26138
rect 19580 26084 19636 26086
rect 19660 26084 19716 26086
rect 19740 26084 19796 26086
rect 19820 26084 19876 26086
rect 19580 25050 19636 25052
rect 19660 25050 19716 25052
rect 19740 25050 19796 25052
rect 19820 25050 19876 25052
rect 19580 24998 19626 25050
rect 19626 24998 19636 25050
rect 19660 24998 19690 25050
rect 19690 24998 19702 25050
rect 19702 24998 19716 25050
rect 19740 24998 19754 25050
rect 19754 24998 19766 25050
rect 19766 24998 19796 25050
rect 19820 24998 19830 25050
rect 19830 24998 19876 25050
rect 19580 24996 19636 24998
rect 19660 24996 19716 24998
rect 19740 24996 19796 24998
rect 19820 24996 19876 24998
rect 19580 23962 19636 23964
rect 19660 23962 19716 23964
rect 19740 23962 19796 23964
rect 19820 23962 19876 23964
rect 19580 23910 19626 23962
rect 19626 23910 19636 23962
rect 19660 23910 19690 23962
rect 19690 23910 19702 23962
rect 19702 23910 19716 23962
rect 19740 23910 19754 23962
rect 19754 23910 19766 23962
rect 19766 23910 19796 23962
rect 19820 23910 19830 23962
rect 19830 23910 19876 23962
rect 19580 23908 19636 23910
rect 19660 23908 19716 23910
rect 19740 23908 19796 23910
rect 19820 23908 19876 23910
rect 19580 22874 19636 22876
rect 19660 22874 19716 22876
rect 19740 22874 19796 22876
rect 19820 22874 19876 22876
rect 19580 22822 19626 22874
rect 19626 22822 19636 22874
rect 19660 22822 19690 22874
rect 19690 22822 19702 22874
rect 19702 22822 19716 22874
rect 19740 22822 19754 22874
rect 19754 22822 19766 22874
rect 19766 22822 19796 22874
rect 19820 22822 19830 22874
rect 19830 22822 19876 22874
rect 19580 22820 19636 22822
rect 19660 22820 19716 22822
rect 19740 22820 19796 22822
rect 19820 22820 19876 22822
rect 19580 21786 19636 21788
rect 19660 21786 19716 21788
rect 19740 21786 19796 21788
rect 19820 21786 19876 21788
rect 19580 21734 19626 21786
rect 19626 21734 19636 21786
rect 19660 21734 19690 21786
rect 19690 21734 19702 21786
rect 19702 21734 19716 21786
rect 19740 21734 19754 21786
rect 19754 21734 19766 21786
rect 19766 21734 19796 21786
rect 19820 21734 19830 21786
rect 19830 21734 19876 21786
rect 19580 21732 19636 21734
rect 19660 21732 19716 21734
rect 19740 21732 19796 21734
rect 19820 21732 19876 21734
rect 19580 20698 19636 20700
rect 19660 20698 19716 20700
rect 19740 20698 19796 20700
rect 19820 20698 19876 20700
rect 19580 20646 19626 20698
rect 19626 20646 19636 20698
rect 19660 20646 19690 20698
rect 19690 20646 19702 20698
rect 19702 20646 19716 20698
rect 19740 20646 19754 20698
rect 19754 20646 19766 20698
rect 19766 20646 19796 20698
rect 19820 20646 19830 20698
rect 19830 20646 19876 20698
rect 19580 20644 19636 20646
rect 19660 20644 19716 20646
rect 19740 20644 19796 20646
rect 19820 20644 19876 20646
rect 19580 19610 19636 19612
rect 19660 19610 19716 19612
rect 19740 19610 19796 19612
rect 19820 19610 19876 19612
rect 19580 19558 19626 19610
rect 19626 19558 19636 19610
rect 19660 19558 19690 19610
rect 19690 19558 19702 19610
rect 19702 19558 19716 19610
rect 19740 19558 19754 19610
rect 19754 19558 19766 19610
rect 19766 19558 19796 19610
rect 19820 19558 19830 19610
rect 19830 19558 19876 19610
rect 19580 19556 19636 19558
rect 19660 19556 19716 19558
rect 19740 19556 19796 19558
rect 19820 19556 19876 19558
rect 19580 18522 19636 18524
rect 19660 18522 19716 18524
rect 19740 18522 19796 18524
rect 19820 18522 19876 18524
rect 19580 18470 19626 18522
rect 19626 18470 19636 18522
rect 19660 18470 19690 18522
rect 19690 18470 19702 18522
rect 19702 18470 19716 18522
rect 19740 18470 19754 18522
rect 19754 18470 19766 18522
rect 19766 18470 19796 18522
rect 19820 18470 19830 18522
rect 19830 18470 19876 18522
rect 19580 18468 19636 18470
rect 19660 18468 19716 18470
rect 19740 18468 19796 18470
rect 19820 18468 19876 18470
rect 19580 17434 19636 17436
rect 19660 17434 19716 17436
rect 19740 17434 19796 17436
rect 19820 17434 19876 17436
rect 19580 17382 19626 17434
rect 19626 17382 19636 17434
rect 19660 17382 19690 17434
rect 19690 17382 19702 17434
rect 19702 17382 19716 17434
rect 19740 17382 19754 17434
rect 19754 17382 19766 17434
rect 19766 17382 19796 17434
rect 19820 17382 19830 17434
rect 19830 17382 19876 17434
rect 19580 17380 19636 17382
rect 19660 17380 19716 17382
rect 19740 17380 19796 17382
rect 19820 17380 19876 17382
rect 19580 16346 19636 16348
rect 19660 16346 19716 16348
rect 19740 16346 19796 16348
rect 19820 16346 19876 16348
rect 19580 16294 19626 16346
rect 19626 16294 19636 16346
rect 19660 16294 19690 16346
rect 19690 16294 19702 16346
rect 19702 16294 19716 16346
rect 19740 16294 19754 16346
rect 19754 16294 19766 16346
rect 19766 16294 19796 16346
rect 19820 16294 19830 16346
rect 19830 16294 19876 16346
rect 19580 16292 19636 16294
rect 19660 16292 19716 16294
rect 19740 16292 19796 16294
rect 19820 16292 19876 16294
rect 19580 15258 19636 15260
rect 19660 15258 19716 15260
rect 19740 15258 19796 15260
rect 19820 15258 19876 15260
rect 19580 15206 19626 15258
rect 19626 15206 19636 15258
rect 19660 15206 19690 15258
rect 19690 15206 19702 15258
rect 19702 15206 19716 15258
rect 19740 15206 19754 15258
rect 19754 15206 19766 15258
rect 19766 15206 19796 15258
rect 19820 15206 19830 15258
rect 19830 15206 19876 15258
rect 19580 15204 19636 15206
rect 19660 15204 19716 15206
rect 19740 15204 19796 15206
rect 19820 15204 19876 15206
rect 19580 14170 19636 14172
rect 19660 14170 19716 14172
rect 19740 14170 19796 14172
rect 19820 14170 19876 14172
rect 19580 14118 19626 14170
rect 19626 14118 19636 14170
rect 19660 14118 19690 14170
rect 19690 14118 19702 14170
rect 19702 14118 19716 14170
rect 19740 14118 19754 14170
rect 19754 14118 19766 14170
rect 19766 14118 19796 14170
rect 19820 14118 19830 14170
rect 19830 14118 19876 14170
rect 19580 14116 19636 14118
rect 19660 14116 19716 14118
rect 19740 14116 19796 14118
rect 19820 14116 19876 14118
rect 19580 13082 19636 13084
rect 19660 13082 19716 13084
rect 19740 13082 19796 13084
rect 19820 13082 19876 13084
rect 19580 13030 19626 13082
rect 19626 13030 19636 13082
rect 19660 13030 19690 13082
rect 19690 13030 19702 13082
rect 19702 13030 19716 13082
rect 19740 13030 19754 13082
rect 19754 13030 19766 13082
rect 19766 13030 19796 13082
rect 19820 13030 19830 13082
rect 19830 13030 19876 13082
rect 19580 13028 19636 13030
rect 19660 13028 19716 13030
rect 19740 13028 19796 13030
rect 19820 13028 19876 13030
rect 19580 11994 19636 11996
rect 19660 11994 19716 11996
rect 19740 11994 19796 11996
rect 19820 11994 19876 11996
rect 19580 11942 19626 11994
rect 19626 11942 19636 11994
rect 19660 11942 19690 11994
rect 19690 11942 19702 11994
rect 19702 11942 19716 11994
rect 19740 11942 19754 11994
rect 19754 11942 19766 11994
rect 19766 11942 19796 11994
rect 19820 11942 19830 11994
rect 19830 11942 19876 11994
rect 19580 11940 19636 11942
rect 19660 11940 19716 11942
rect 19740 11940 19796 11942
rect 19820 11940 19876 11942
rect 19580 10906 19636 10908
rect 19660 10906 19716 10908
rect 19740 10906 19796 10908
rect 19820 10906 19876 10908
rect 19580 10854 19626 10906
rect 19626 10854 19636 10906
rect 19660 10854 19690 10906
rect 19690 10854 19702 10906
rect 19702 10854 19716 10906
rect 19740 10854 19754 10906
rect 19754 10854 19766 10906
rect 19766 10854 19796 10906
rect 19820 10854 19830 10906
rect 19830 10854 19876 10906
rect 19580 10852 19636 10854
rect 19660 10852 19716 10854
rect 19740 10852 19796 10854
rect 19820 10852 19876 10854
rect 19580 9818 19636 9820
rect 19660 9818 19716 9820
rect 19740 9818 19796 9820
rect 19820 9818 19876 9820
rect 19580 9766 19626 9818
rect 19626 9766 19636 9818
rect 19660 9766 19690 9818
rect 19690 9766 19702 9818
rect 19702 9766 19716 9818
rect 19740 9766 19754 9818
rect 19754 9766 19766 9818
rect 19766 9766 19796 9818
rect 19820 9766 19830 9818
rect 19830 9766 19876 9818
rect 19580 9764 19636 9766
rect 19660 9764 19716 9766
rect 19740 9764 19796 9766
rect 19820 9764 19876 9766
rect 19580 8730 19636 8732
rect 19660 8730 19716 8732
rect 19740 8730 19796 8732
rect 19820 8730 19876 8732
rect 19580 8678 19626 8730
rect 19626 8678 19636 8730
rect 19660 8678 19690 8730
rect 19690 8678 19702 8730
rect 19702 8678 19716 8730
rect 19740 8678 19754 8730
rect 19754 8678 19766 8730
rect 19766 8678 19796 8730
rect 19820 8678 19830 8730
rect 19830 8678 19876 8730
rect 19580 8676 19636 8678
rect 19660 8676 19716 8678
rect 19740 8676 19796 8678
rect 19820 8676 19876 8678
rect 19580 7642 19636 7644
rect 19660 7642 19716 7644
rect 19740 7642 19796 7644
rect 19820 7642 19876 7644
rect 19580 7590 19626 7642
rect 19626 7590 19636 7642
rect 19660 7590 19690 7642
rect 19690 7590 19702 7642
rect 19702 7590 19716 7642
rect 19740 7590 19754 7642
rect 19754 7590 19766 7642
rect 19766 7590 19796 7642
rect 19820 7590 19830 7642
rect 19830 7590 19876 7642
rect 19580 7588 19636 7590
rect 19660 7588 19716 7590
rect 19740 7588 19796 7590
rect 19820 7588 19876 7590
rect 19580 6554 19636 6556
rect 19660 6554 19716 6556
rect 19740 6554 19796 6556
rect 19820 6554 19876 6556
rect 19580 6502 19626 6554
rect 19626 6502 19636 6554
rect 19660 6502 19690 6554
rect 19690 6502 19702 6554
rect 19702 6502 19716 6554
rect 19740 6502 19754 6554
rect 19754 6502 19766 6554
rect 19766 6502 19796 6554
rect 19820 6502 19830 6554
rect 19830 6502 19876 6554
rect 19580 6500 19636 6502
rect 19660 6500 19716 6502
rect 19740 6500 19796 6502
rect 19820 6500 19876 6502
rect 19580 5466 19636 5468
rect 19660 5466 19716 5468
rect 19740 5466 19796 5468
rect 19820 5466 19876 5468
rect 19580 5414 19626 5466
rect 19626 5414 19636 5466
rect 19660 5414 19690 5466
rect 19690 5414 19702 5466
rect 19702 5414 19716 5466
rect 19740 5414 19754 5466
rect 19754 5414 19766 5466
rect 19766 5414 19796 5466
rect 19820 5414 19830 5466
rect 19830 5414 19876 5466
rect 19580 5412 19636 5414
rect 19660 5412 19716 5414
rect 19740 5412 19796 5414
rect 19820 5412 19876 5414
rect 19580 4378 19636 4380
rect 19660 4378 19716 4380
rect 19740 4378 19796 4380
rect 19820 4378 19876 4380
rect 19580 4326 19626 4378
rect 19626 4326 19636 4378
rect 19660 4326 19690 4378
rect 19690 4326 19702 4378
rect 19702 4326 19716 4378
rect 19740 4326 19754 4378
rect 19754 4326 19766 4378
rect 19766 4326 19796 4378
rect 19820 4326 19830 4378
rect 19830 4326 19876 4378
rect 19580 4324 19636 4326
rect 19660 4324 19716 4326
rect 19740 4324 19796 4326
rect 19820 4324 19876 4326
rect 19580 3290 19636 3292
rect 19660 3290 19716 3292
rect 19740 3290 19796 3292
rect 19820 3290 19876 3292
rect 19580 3238 19626 3290
rect 19626 3238 19636 3290
rect 19660 3238 19690 3290
rect 19690 3238 19702 3290
rect 19702 3238 19716 3290
rect 19740 3238 19754 3290
rect 19754 3238 19766 3290
rect 19766 3238 19796 3290
rect 19820 3238 19830 3290
rect 19830 3238 19876 3290
rect 19580 3236 19636 3238
rect 19660 3236 19716 3238
rect 19740 3236 19796 3238
rect 19820 3236 19876 3238
rect 34940 59322 34996 59324
rect 35020 59322 35076 59324
rect 35100 59322 35156 59324
rect 35180 59322 35236 59324
rect 34940 59270 34986 59322
rect 34986 59270 34996 59322
rect 35020 59270 35050 59322
rect 35050 59270 35062 59322
rect 35062 59270 35076 59322
rect 35100 59270 35114 59322
rect 35114 59270 35126 59322
rect 35126 59270 35156 59322
rect 35180 59270 35190 59322
rect 35190 59270 35236 59322
rect 34940 59268 34996 59270
rect 35020 59268 35076 59270
rect 35100 59268 35156 59270
rect 35180 59268 35236 59270
rect 34940 58234 34996 58236
rect 35020 58234 35076 58236
rect 35100 58234 35156 58236
rect 35180 58234 35236 58236
rect 34940 58182 34986 58234
rect 34986 58182 34996 58234
rect 35020 58182 35050 58234
rect 35050 58182 35062 58234
rect 35062 58182 35076 58234
rect 35100 58182 35114 58234
rect 35114 58182 35126 58234
rect 35126 58182 35156 58234
rect 35180 58182 35190 58234
rect 35190 58182 35236 58234
rect 34940 58180 34996 58182
rect 35020 58180 35076 58182
rect 35100 58180 35156 58182
rect 35180 58180 35236 58182
rect 34940 57146 34996 57148
rect 35020 57146 35076 57148
rect 35100 57146 35156 57148
rect 35180 57146 35236 57148
rect 34940 57094 34986 57146
rect 34986 57094 34996 57146
rect 35020 57094 35050 57146
rect 35050 57094 35062 57146
rect 35062 57094 35076 57146
rect 35100 57094 35114 57146
rect 35114 57094 35126 57146
rect 35126 57094 35156 57146
rect 35180 57094 35190 57146
rect 35190 57094 35236 57146
rect 34940 57092 34996 57094
rect 35020 57092 35076 57094
rect 35100 57092 35156 57094
rect 35180 57092 35236 57094
rect 34940 56058 34996 56060
rect 35020 56058 35076 56060
rect 35100 56058 35156 56060
rect 35180 56058 35236 56060
rect 34940 56006 34986 56058
rect 34986 56006 34996 56058
rect 35020 56006 35050 56058
rect 35050 56006 35062 56058
rect 35062 56006 35076 56058
rect 35100 56006 35114 56058
rect 35114 56006 35126 56058
rect 35126 56006 35156 56058
rect 35180 56006 35190 56058
rect 35190 56006 35236 56058
rect 34940 56004 34996 56006
rect 35020 56004 35076 56006
rect 35100 56004 35156 56006
rect 35180 56004 35236 56006
rect 34940 54970 34996 54972
rect 35020 54970 35076 54972
rect 35100 54970 35156 54972
rect 35180 54970 35236 54972
rect 34940 54918 34986 54970
rect 34986 54918 34996 54970
rect 35020 54918 35050 54970
rect 35050 54918 35062 54970
rect 35062 54918 35076 54970
rect 35100 54918 35114 54970
rect 35114 54918 35126 54970
rect 35126 54918 35156 54970
rect 35180 54918 35190 54970
rect 35190 54918 35236 54970
rect 34940 54916 34996 54918
rect 35020 54916 35076 54918
rect 35100 54916 35156 54918
rect 35180 54916 35236 54918
rect 34940 53882 34996 53884
rect 35020 53882 35076 53884
rect 35100 53882 35156 53884
rect 35180 53882 35236 53884
rect 34940 53830 34986 53882
rect 34986 53830 34996 53882
rect 35020 53830 35050 53882
rect 35050 53830 35062 53882
rect 35062 53830 35076 53882
rect 35100 53830 35114 53882
rect 35114 53830 35126 53882
rect 35126 53830 35156 53882
rect 35180 53830 35190 53882
rect 35190 53830 35236 53882
rect 34940 53828 34996 53830
rect 35020 53828 35076 53830
rect 35100 53828 35156 53830
rect 35180 53828 35236 53830
rect 34940 52794 34996 52796
rect 35020 52794 35076 52796
rect 35100 52794 35156 52796
rect 35180 52794 35236 52796
rect 34940 52742 34986 52794
rect 34986 52742 34996 52794
rect 35020 52742 35050 52794
rect 35050 52742 35062 52794
rect 35062 52742 35076 52794
rect 35100 52742 35114 52794
rect 35114 52742 35126 52794
rect 35126 52742 35156 52794
rect 35180 52742 35190 52794
rect 35190 52742 35236 52794
rect 34940 52740 34996 52742
rect 35020 52740 35076 52742
rect 35100 52740 35156 52742
rect 35180 52740 35236 52742
rect 34940 51706 34996 51708
rect 35020 51706 35076 51708
rect 35100 51706 35156 51708
rect 35180 51706 35236 51708
rect 34940 51654 34986 51706
rect 34986 51654 34996 51706
rect 35020 51654 35050 51706
rect 35050 51654 35062 51706
rect 35062 51654 35076 51706
rect 35100 51654 35114 51706
rect 35114 51654 35126 51706
rect 35126 51654 35156 51706
rect 35180 51654 35190 51706
rect 35190 51654 35236 51706
rect 34940 51652 34996 51654
rect 35020 51652 35076 51654
rect 35100 51652 35156 51654
rect 35180 51652 35236 51654
rect 34940 50618 34996 50620
rect 35020 50618 35076 50620
rect 35100 50618 35156 50620
rect 35180 50618 35236 50620
rect 34940 50566 34986 50618
rect 34986 50566 34996 50618
rect 35020 50566 35050 50618
rect 35050 50566 35062 50618
rect 35062 50566 35076 50618
rect 35100 50566 35114 50618
rect 35114 50566 35126 50618
rect 35126 50566 35156 50618
rect 35180 50566 35190 50618
rect 35190 50566 35236 50618
rect 34940 50564 34996 50566
rect 35020 50564 35076 50566
rect 35100 50564 35156 50566
rect 35180 50564 35236 50566
rect 34940 49530 34996 49532
rect 35020 49530 35076 49532
rect 35100 49530 35156 49532
rect 35180 49530 35236 49532
rect 34940 49478 34986 49530
rect 34986 49478 34996 49530
rect 35020 49478 35050 49530
rect 35050 49478 35062 49530
rect 35062 49478 35076 49530
rect 35100 49478 35114 49530
rect 35114 49478 35126 49530
rect 35126 49478 35156 49530
rect 35180 49478 35190 49530
rect 35190 49478 35236 49530
rect 34940 49476 34996 49478
rect 35020 49476 35076 49478
rect 35100 49476 35156 49478
rect 35180 49476 35236 49478
rect 34940 48442 34996 48444
rect 35020 48442 35076 48444
rect 35100 48442 35156 48444
rect 35180 48442 35236 48444
rect 34940 48390 34986 48442
rect 34986 48390 34996 48442
rect 35020 48390 35050 48442
rect 35050 48390 35062 48442
rect 35062 48390 35076 48442
rect 35100 48390 35114 48442
rect 35114 48390 35126 48442
rect 35126 48390 35156 48442
rect 35180 48390 35190 48442
rect 35190 48390 35236 48442
rect 34940 48388 34996 48390
rect 35020 48388 35076 48390
rect 35100 48388 35156 48390
rect 35180 48388 35236 48390
rect 34940 47354 34996 47356
rect 35020 47354 35076 47356
rect 35100 47354 35156 47356
rect 35180 47354 35236 47356
rect 34940 47302 34986 47354
rect 34986 47302 34996 47354
rect 35020 47302 35050 47354
rect 35050 47302 35062 47354
rect 35062 47302 35076 47354
rect 35100 47302 35114 47354
rect 35114 47302 35126 47354
rect 35126 47302 35156 47354
rect 35180 47302 35190 47354
rect 35190 47302 35236 47354
rect 34940 47300 34996 47302
rect 35020 47300 35076 47302
rect 35100 47300 35156 47302
rect 35180 47300 35236 47302
rect 34940 46266 34996 46268
rect 35020 46266 35076 46268
rect 35100 46266 35156 46268
rect 35180 46266 35236 46268
rect 34940 46214 34986 46266
rect 34986 46214 34996 46266
rect 35020 46214 35050 46266
rect 35050 46214 35062 46266
rect 35062 46214 35076 46266
rect 35100 46214 35114 46266
rect 35114 46214 35126 46266
rect 35126 46214 35156 46266
rect 35180 46214 35190 46266
rect 35190 46214 35236 46266
rect 34940 46212 34996 46214
rect 35020 46212 35076 46214
rect 35100 46212 35156 46214
rect 35180 46212 35236 46214
rect 34940 45178 34996 45180
rect 35020 45178 35076 45180
rect 35100 45178 35156 45180
rect 35180 45178 35236 45180
rect 34940 45126 34986 45178
rect 34986 45126 34996 45178
rect 35020 45126 35050 45178
rect 35050 45126 35062 45178
rect 35062 45126 35076 45178
rect 35100 45126 35114 45178
rect 35114 45126 35126 45178
rect 35126 45126 35156 45178
rect 35180 45126 35190 45178
rect 35190 45126 35236 45178
rect 34940 45124 34996 45126
rect 35020 45124 35076 45126
rect 35100 45124 35156 45126
rect 35180 45124 35236 45126
rect 34940 44090 34996 44092
rect 35020 44090 35076 44092
rect 35100 44090 35156 44092
rect 35180 44090 35236 44092
rect 34940 44038 34986 44090
rect 34986 44038 34996 44090
rect 35020 44038 35050 44090
rect 35050 44038 35062 44090
rect 35062 44038 35076 44090
rect 35100 44038 35114 44090
rect 35114 44038 35126 44090
rect 35126 44038 35156 44090
rect 35180 44038 35190 44090
rect 35190 44038 35236 44090
rect 34940 44036 34996 44038
rect 35020 44036 35076 44038
rect 35100 44036 35156 44038
rect 35180 44036 35236 44038
rect 34940 43002 34996 43004
rect 35020 43002 35076 43004
rect 35100 43002 35156 43004
rect 35180 43002 35236 43004
rect 34940 42950 34986 43002
rect 34986 42950 34996 43002
rect 35020 42950 35050 43002
rect 35050 42950 35062 43002
rect 35062 42950 35076 43002
rect 35100 42950 35114 43002
rect 35114 42950 35126 43002
rect 35126 42950 35156 43002
rect 35180 42950 35190 43002
rect 35190 42950 35236 43002
rect 34940 42948 34996 42950
rect 35020 42948 35076 42950
rect 35100 42948 35156 42950
rect 35180 42948 35236 42950
rect 34940 41914 34996 41916
rect 35020 41914 35076 41916
rect 35100 41914 35156 41916
rect 35180 41914 35236 41916
rect 34940 41862 34986 41914
rect 34986 41862 34996 41914
rect 35020 41862 35050 41914
rect 35050 41862 35062 41914
rect 35062 41862 35076 41914
rect 35100 41862 35114 41914
rect 35114 41862 35126 41914
rect 35126 41862 35156 41914
rect 35180 41862 35190 41914
rect 35190 41862 35236 41914
rect 34940 41860 34996 41862
rect 35020 41860 35076 41862
rect 35100 41860 35156 41862
rect 35180 41860 35236 41862
rect 34940 40826 34996 40828
rect 35020 40826 35076 40828
rect 35100 40826 35156 40828
rect 35180 40826 35236 40828
rect 34940 40774 34986 40826
rect 34986 40774 34996 40826
rect 35020 40774 35050 40826
rect 35050 40774 35062 40826
rect 35062 40774 35076 40826
rect 35100 40774 35114 40826
rect 35114 40774 35126 40826
rect 35126 40774 35156 40826
rect 35180 40774 35190 40826
rect 35190 40774 35236 40826
rect 34940 40772 34996 40774
rect 35020 40772 35076 40774
rect 35100 40772 35156 40774
rect 35180 40772 35236 40774
rect 34940 39738 34996 39740
rect 35020 39738 35076 39740
rect 35100 39738 35156 39740
rect 35180 39738 35236 39740
rect 34940 39686 34986 39738
rect 34986 39686 34996 39738
rect 35020 39686 35050 39738
rect 35050 39686 35062 39738
rect 35062 39686 35076 39738
rect 35100 39686 35114 39738
rect 35114 39686 35126 39738
rect 35126 39686 35156 39738
rect 35180 39686 35190 39738
rect 35190 39686 35236 39738
rect 34940 39684 34996 39686
rect 35020 39684 35076 39686
rect 35100 39684 35156 39686
rect 35180 39684 35236 39686
rect 34940 38650 34996 38652
rect 35020 38650 35076 38652
rect 35100 38650 35156 38652
rect 35180 38650 35236 38652
rect 34940 38598 34986 38650
rect 34986 38598 34996 38650
rect 35020 38598 35050 38650
rect 35050 38598 35062 38650
rect 35062 38598 35076 38650
rect 35100 38598 35114 38650
rect 35114 38598 35126 38650
rect 35126 38598 35156 38650
rect 35180 38598 35190 38650
rect 35190 38598 35236 38650
rect 34940 38596 34996 38598
rect 35020 38596 35076 38598
rect 35100 38596 35156 38598
rect 35180 38596 35236 38598
rect 34940 37562 34996 37564
rect 35020 37562 35076 37564
rect 35100 37562 35156 37564
rect 35180 37562 35236 37564
rect 34940 37510 34986 37562
rect 34986 37510 34996 37562
rect 35020 37510 35050 37562
rect 35050 37510 35062 37562
rect 35062 37510 35076 37562
rect 35100 37510 35114 37562
rect 35114 37510 35126 37562
rect 35126 37510 35156 37562
rect 35180 37510 35190 37562
rect 35190 37510 35236 37562
rect 34940 37508 34996 37510
rect 35020 37508 35076 37510
rect 35100 37508 35156 37510
rect 35180 37508 35236 37510
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
rect 19580 2202 19636 2204
rect 19660 2202 19716 2204
rect 19740 2202 19796 2204
rect 19820 2202 19876 2204
rect 19580 2150 19626 2202
rect 19626 2150 19636 2202
rect 19660 2150 19690 2202
rect 19690 2150 19702 2202
rect 19702 2150 19716 2202
rect 19740 2150 19754 2202
rect 19754 2150 19766 2202
rect 19766 2150 19796 2202
rect 19820 2150 19830 2202
rect 19830 2150 19876 2202
rect 19580 2148 19636 2150
rect 19660 2148 19716 2150
rect 19740 2148 19796 2150
rect 19820 2148 19876 2150
rect 50300 117530 50356 117532
rect 50380 117530 50436 117532
rect 50460 117530 50516 117532
rect 50540 117530 50596 117532
rect 50300 117478 50346 117530
rect 50346 117478 50356 117530
rect 50380 117478 50410 117530
rect 50410 117478 50422 117530
rect 50422 117478 50436 117530
rect 50460 117478 50474 117530
rect 50474 117478 50486 117530
rect 50486 117478 50516 117530
rect 50540 117478 50550 117530
rect 50550 117478 50596 117530
rect 50300 117476 50356 117478
rect 50380 117476 50436 117478
rect 50460 117476 50516 117478
rect 50540 117476 50596 117478
rect 50300 116442 50356 116444
rect 50380 116442 50436 116444
rect 50460 116442 50516 116444
rect 50540 116442 50596 116444
rect 50300 116390 50346 116442
rect 50346 116390 50356 116442
rect 50380 116390 50410 116442
rect 50410 116390 50422 116442
rect 50422 116390 50436 116442
rect 50460 116390 50474 116442
rect 50474 116390 50486 116442
rect 50486 116390 50516 116442
rect 50540 116390 50550 116442
rect 50550 116390 50596 116442
rect 50300 116388 50356 116390
rect 50380 116388 50436 116390
rect 50460 116388 50516 116390
rect 50540 116388 50596 116390
rect 50300 115354 50356 115356
rect 50380 115354 50436 115356
rect 50460 115354 50516 115356
rect 50540 115354 50596 115356
rect 50300 115302 50346 115354
rect 50346 115302 50356 115354
rect 50380 115302 50410 115354
rect 50410 115302 50422 115354
rect 50422 115302 50436 115354
rect 50460 115302 50474 115354
rect 50474 115302 50486 115354
rect 50486 115302 50516 115354
rect 50540 115302 50550 115354
rect 50550 115302 50596 115354
rect 50300 115300 50356 115302
rect 50380 115300 50436 115302
rect 50460 115300 50516 115302
rect 50540 115300 50596 115302
rect 50300 114266 50356 114268
rect 50380 114266 50436 114268
rect 50460 114266 50516 114268
rect 50540 114266 50596 114268
rect 50300 114214 50346 114266
rect 50346 114214 50356 114266
rect 50380 114214 50410 114266
rect 50410 114214 50422 114266
rect 50422 114214 50436 114266
rect 50460 114214 50474 114266
rect 50474 114214 50486 114266
rect 50486 114214 50516 114266
rect 50540 114214 50550 114266
rect 50550 114214 50596 114266
rect 50300 114212 50356 114214
rect 50380 114212 50436 114214
rect 50460 114212 50516 114214
rect 50540 114212 50596 114214
rect 50300 113178 50356 113180
rect 50380 113178 50436 113180
rect 50460 113178 50516 113180
rect 50540 113178 50596 113180
rect 50300 113126 50346 113178
rect 50346 113126 50356 113178
rect 50380 113126 50410 113178
rect 50410 113126 50422 113178
rect 50422 113126 50436 113178
rect 50460 113126 50474 113178
rect 50474 113126 50486 113178
rect 50486 113126 50516 113178
rect 50540 113126 50550 113178
rect 50550 113126 50596 113178
rect 50300 113124 50356 113126
rect 50380 113124 50436 113126
rect 50460 113124 50516 113126
rect 50540 113124 50596 113126
rect 50300 112090 50356 112092
rect 50380 112090 50436 112092
rect 50460 112090 50516 112092
rect 50540 112090 50596 112092
rect 50300 112038 50346 112090
rect 50346 112038 50356 112090
rect 50380 112038 50410 112090
rect 50410 112038 50422 112090
rect 50422 112038 50436 112090
rect 50460 112038 50474 112090
rect 50474 112038 50486 112090
rect 50486 112038 50516 112090
rect 50540 112038 50550 112090
rect 50550 112038 50596 112090
rect 50300 112036 50356 112038
rect 50380 112036 50436 112038
rect 50460 112036 50516 112038
rect 50540 112036 50596 112038
rect 50300 111002 50356 111004
rect 50380 111002 50436 111004
rect 50460 111002 50516 111004
rect 50540 111002 50596 111004
rect 50300 110950 50346 111002
rect 50346 110950 50356 111002
rect 50380 110950 50410 111002
rect 50410 110950 50422 111002
rect 50422 110950 50436 111002
rect 50460 110950 50474 111002
rect 50474 110950 50486 111002
rect 50486 110950 50516 111002
rect 50540 110950 50550 111002
rect 50550 110950 50596 111002
rect 50300 110948 50356 110950
rect 50380 110948 50436 110950
rect 50460 110948 50516 110950
rect 50540 110948 50596 110950
rect 50300 109914 50356 109916
rect 50380 109914 50436 109916
rect 50460 109914 50516 109916
rect 50540 109914 50596 109916
rect 50300 109862 50346 109914
rect 50346 109862 50356 109914
rect 50380 109862 50410 109914
rect 50410 109862 50422 109914
rect 50422 109862 50436 109914
rect 50460 109862 50474 109914
rect 50474 109862 50486 109914
rect 50486 109862 50516 109914
rect 50540 109862 50550 109914
rect 50550 109862 50596 109914
rect 50300 109860 50356 109862
rect 50380 109860 50436 109862
rect 50460 109860 50516 109862
rect 50540 109860 50596 109862
rect 50300 108826 50356 108828
rect 50380 108826 50436 108828
rect 50460 108826 50516 108828
rect 50540 108826 50596 108828
rect 50300 108774 50346 108826
rect 50346 108774 50356 108826
rect 50380 108774 50410 108826
rect 50410 108774 50422 108826
rect 50422 108774 50436 108826
rect 50460 108774 50474 108826
rect 50474 108774 50486 108826
rect 50486 108774 50516 108826
rect 50540 108774 50550 108826
rect 50550 108774 50596 108826
rect 50300 108772 50356 108774
rect 50380 108772 50436 108774
rect 50460 108772 50516 108774
rect 50540 108772 50596 108774
rect 50300 107738 50356 107740
rect 50380 107738 50436 107740
rect 50460 107738 50516 107740
rect 50540 107738 50596 107740
rect 50300 107686 50346 107738
rect 50346 107686 50356 107738
rect 50380 107686 50410 107738
rect 50410 107686 50422 107738
rect 50422 107686 50436 107738
rect 50460 107686 50474 107738
rect 50474 107686 50486 107738
rect 50486 107686 50516 107738
rect 50540 107686 50550 107738
rect 50550 107686 50596 107738
rect 50300 107684 50356 107686
rect 50380 107684 50436 107686
rect 50460 107684 50516 107686
rect 50540 107684 50596 107686
rect 50300 106650 50356 106652
rect 50380 106650 50436 106652
rect 50460 106650 50516 106652
rect 50540 106650 50596 106652
rect 50300 106598 50346 106650
rect 50346 106598 50356 106650
rect 50380 106598 50410 106650
rect 50410 106598 50422 106650
rect 50422 106598 50436 106650
rect 50460 106598 50474 106650
rect 50474 106598 50486 106650
rect 50486 106598 50516 106650
rect 50540 106598 50550 106650
rect 50550 106598 50596 106650
rect 50300 106596 50356 106598
rect 50380 106596 50436 106598
rect 50460 106596 50516 106598
rect 50540 106596 50596 106598
rect 50300 105562 50356 105564
rect 50380 105562 50436 105564
rect 50460 105562 50516 105564
rect 50540 105562 50596 105564
rect 50300 105510 50346 105562
rect 50346 105510 50356 105562
rect 50380 105510 50410 105562
rect 50410 105510 50422 105562
rect 50422 105510 50436 105562
rect 50460 105510 50474 105562
rect 50474 105510 50486 105562
rect 50486 105510 50516 105562
rect 50540 105510 50550 105562
rect 50550 105510 50596 105562
rect 50300 105508 50356 105510
rect 50380 105508 50436 105510
rect 50460 105508 50516 105510
rect 50540 105508 50596 105510
rect 50300 104474 50356 104476
rect 50380 104474 50436 104476
rect 50460 104474 50516 104476
rect 50540 104474 50596 104476
rect 50300 104422 50346 104474
rect 50346 104422 50356 104474
rect 50380 104422 50410 104474
rect 50410 104422 50422 104474
rect 50422 104422 50436 104474
rect 50460 104422 50474 104474
rect 50474 104422 50486 104474
rect 50486 104422 50516 104474
rect 50540 104422 50550 104474
rect 50550 104422 50596 104474
rect 50300 104420 50356 104422
rect 50380 104420 50436 104422
rect 50460 104420 50516 104422
rect 50540 104420 50596 104422
rect 50300 103386 50356 103388
rect 50380 103386 50436 103388
rect 50460 103386 50516 103388
rect 50540 103386 50596 103388
rect 50300 103334 50346 103386
rect 50346 103334 50356 103386
rect 50380 103334 50410 103386
rect 50410 103334 50422 103386
rect 50422 103334 50436 103386
rect 50460 103334 50474 103386
rect 50474 103334 50486 103386
rect 50486 103334 50516 103386
rect 50540 103334 50550 103386
rect 50550 103334 50596 103386
rect 50300 103332 50356 103334
rect 50380 103332 50436 103334
rect 50460 103332 50516 103334
rect 50540 103332 50596 103334
rect 50300 102298 50356 102300
rect 50380 102298 50436 102300
rect 50460 102298 50516 102300
rect 50540 102298 50596 102300
rect 50300 102246 50346 102298
rect 50346 102246 50356 102298
rect 50380 102246 50410 102298
rect 50410 102246 50422 102298
rect 50422 102246 50436 102298
rect 50460 102246 50474 102298
rect 50474 102246 50486 102298
rect 50486 102246 50516 102298
rect 50540 102246 50550 102298
rect 50550 102246 50596 102298
rect 50300 102244 50356 102246
rect 50380 102244 50436 102246
rect 50460 102244 50516 102246
rect 50540 102244 50596 102246
rect 50300 101210 50356 101212
rect 50380 101210 50436 101212
rect 50460 101210 50516 101212
rect 50540 101210 50596 101212
rect 50300 101158 50346 101210
rect 50346 101158 50356 101210
rect 50380 101158 50410 101210
rect 50410 101158 50422 101210
rect 50422 101158 50436 101210
rect 50460 101158 50474 101210
rect 50474 101158 50486 101210
rect 50486 101158 50516 101210
rect 50540 101158 50550 101210
rect 50550 101158 50596 101210
rect 50300 101156 50356 101158
rect 50380 101156 50436 101158
rect 50460 101156 50516 101158
rect 50540 101156 50596 101158
rect 50300 100122 50356 100124
rect 50380 100122 50436 100124
rect 50460 100122 50516 100124
rect 50540 100122 50596 100124
rect 50300 100070 50346 100122
rect 50346 100070 50356 100122
rect 50380 100070 50410 100122
rect 50410 100070 50422 100122
rect 50422 100070 50436 100122
rect 50460 100070 50474 100122
rect 50474 100070 50486 100122
rect 50486 100070 50516 100122
rect 50540 100070 50550 100122
rect 50550 100070 50596 100122
rect 50300 100068 50356 100070
rect 50380 100068 50436 100070
rect 50460 100068 50516 100070
rect 50540 100068 50596 100070
rect 50300 99034 50356 99036
rect 50380 99034 50436 99036
rect 50460 99034 50516 99036
rect 50540 99034 50596 99036
rect 50300 98982 50346 99034
rect 50346 98982 50356 99034
rect 50380 98982 50410 99034
rect 50410 98982 50422 99034
rect 50422 98982 50436 99034
rect 50460 98982 50474 99034
rect 50474 98982 50486 99034
rect 50486 98982 50516 99034
rect 50540 98982 50550 99034
rect 50550 98982 50596 99034
rect 50300 98980 50356 98982
rect 50380 98980 50436 98982
rect 50460 98980 50516 98982
rect 50540 98980 50596 98982
rect 50300 97946 50356 97948
rect 50380 97946 50436 97948
rect 50460 97946 50516 97948
rect 50540 97946 50596 97948
rect 50300 97894 50346 97946
rect 50346 97894 50356 97946
rect 50380 97894 50410 97946
rect 50410 97894 50422 97946
rect 50422 97894 50436 97946
rect 50460 97894 50474 97946
rect 50474 97894 50486 97946
rect 50486 97894 50516 97946
rect 50540 97894 50550 97946
rect 50550 97894 50596 97946
rect 50300 97892 50356 97894
rect 50380 97892 50436 97894
rect 50460 97892 50516 97894
rect 50540 97892 50596 97894
rect 50300 96858 50356 96860
rect 50380 96858 50436 96860
rect 50460 96858 50516 96860
rect 50540 96858 50596 96860
rect 50300 96806 50346 96858
rect 50346 96806 50356 96858
rect 50380 96806 50410 96858
rect 50410 96806 50422 96858
rect 50422 96806 50436 96858
rect 50460 96806 50474 96858
rect 50474 96806 50486 96858
rect 50486 96806 50516 96858
rect 50540 96806 50550 96858
rect 50550 96806 50596 96858
rect 50300 96804 50356 96806
rect 50380 96804 50436 96806
rect 50460 96804 50516 96806
rect 50540 96804 50596 96806
rect 50300 95770 50356 95772
rect 50380 95770 50436 95772
rect 50460 95770 50516 95772
rect 50540 95770 50596 95772
rect 50300 95718 50346 95770
rect 50346 95718 50356 95770
rect 50380 95718 50410 95770
rect 50410 95718 50422 95770
rect 50422 95718 50436 95770
rect 50460 95718 50474 95770
rect 50474 95718 50486 95770
rect 50486 95718 50516 95770
rect 50540 95718 50550 95770
rect 50550 95718 50596 95770
rect 50300 95716 50356 95718
rect 50380 95716 50436 95718
rect 50460 95716 50516 95718
rect 50540 95716 50596 95718
rect 50300 94682 50356 94684
rect 50380 94682 50436 94684
rect 50460 94682 50516 94684
rect 50540 94682 50596 94684
rect 50300 94630 50346 94682
rect 50346 94630 50356 94682
rect 50380 94630 50410 94682
rect 50410 94630 50422 94682
rect 50422 94630 50436 94682
rect 50460 94630 50474 94682
rect 50474 94630 50486 94682
rect 50486 94630 50516 94682
rect 50540 94630 50550 94682
rect 50550 94630 50596 94682
rect 50300 94628 50356 94630
rect 50380 94628 50436 94630
rect 50460 94628 50516 94630
rect 50540 94628 50596 94630
rect 50300 93594 50356 93596
rect 50380 93594 50436 93596
rect 50460 93594 50516 93596
rect 50540 93594 50596 93596
rect 50300 93542 50346 93594
rect 50346 93542 50356 93594
rect 50380 93542 50410 93594
rect 50410 93542 50422 93594
rect 50422 93542 50436 93594
rect 50460 93542 50474 93594
rect 50474 93542 50486 93594
rect 50486 93542 50516 93594
rect 50540 93542 50550 93594
rect 50550 93542 50596 93594
rect 50300 93540 50356 93542
rect 50380 93540 50436 93542
rect 50460 93540 50516 93542
rect 50540 93540 50596 93542
rect 50300 92506 50356 92508
rect 50380 92506 50436 92508
rect 50460 92506 50516 92508
rect 50540 92506 50596 92508
rect 50300 92454 50346 92506
rect 50346 92454 50356 92506
rect 50380 92454 50410 92506
rect 50410 92454 50422 92506
rect 50422 92454 50436 92506
rect 50460 92454 50474 92506
rect 50474 92454 50486 92506
rect 50486 92454 50516 92506
rect 50540 92454 50550 92506
rect 50550 92454 50596 92506
rect 50300 92452 50356 92454
rect 50380 92452 50436 92454
rect 50460 92452 50516 92454
rect 50540 92452 50596 92454
rect 50300 91418 50356 91420
rect 50380 91418 50436 91420
rect 50460 91418 50516 91420
rect 50540 91418 50596 91420
rect 50300 91366 50346 91418
rect 50346 91366 50356 91418
rect 50380 91366 50410 91418
rect 50410 91366 50422 91418
rect 50422 91366 50436 91418
rect 50460 91366 50474 91418
rect 50474 91366 50486 91418
rect 50486 91366 50516 91418
rect 50540 91366 50550 91418
rect 50550 91366 50596 91418
rect 50300 91364 50356 91366
rect 50380 91364 50436 91366
rect 50460 91364 50516 91366
rect 50540 91364 50596 91366
rect 50300 90330 50356 90332
rect 50380 90330 50436 90332
rect 50460 90330 50516 90332
rect 50540 90330 50596 90332
rect 50300 90278 50346 90330
rect 50346 90278 50356 90330
rect 50380 90278 50410 90330
rect 50410 90278 50422 90330
rect 50422 90278 50436 90330
rect 50460 90278 50474 90330
rect 50474 90278 50486 90330
rect 50486 90278 50516 90330
rect 50540 90278 50550 90330
rect 50550 90278 50596 90330
rect 50300 90276 50356 90278
rect 50380 90276 50436 90278
rect 50460 90276 50516 90278
rect 50540 90276 50596 90278
rect 50300 89242 50356 89244
rect 50380 89242 50436 89244
rect 50460 89242 50516 89244
rect 50540 89242 50596 89244
rect 50300 89190 50346 89242
rect 50346 89190 50356 89242
rect 50380 89190 50410 89242
rect 50410 89190 50422 89242
rect 50422 89190 50436 89242
rect 50460 89190 50474 89242
rect 50474 89190 50486 89242
rect 50486 89190 50516 89242
rect 50540 89190 50550 89242
rect 50550 89190 50596 89242
rect 50300 89188 50356 89190
rect 50380 89188 50436 89190
rect 50460 89188 50516 89190
rect 50540 89188 50596 89190
rect 50300 88154 50356 88156
rect 50380 88154 50436 88156
rect 50460 88154 50516 88156
rect 50540 88154 50596 88156
rect 50300 88102 50346 88154
rect 50346 88102 50356 88154
rect 50380 88102 50410 88154
rect 50410 88102 50422 88154
rect 50422 88102 50436 88154
rect 50460 88102 50474 88154
rect 50474 88102 50486 88154
rect 50486 88102 50516 88154
rect 50540 88102 50550 88154
rect 50550 88102 50596 88154
rect 50300 88100 50356 88102
rect 50380 88100 50436 88102
rect 50460 88100 50516 88102
rect 50540 88100 50596 88102
rect 50300 87066 50356 87068
rect 50380 87066 50436 87068
rect 50460 87066 50516 87068
rect 50540 87066 50596 87068
rect 50300 87014 50346 87066
rect 50346 87014 50356 87066
rect 50380 87014 50410 87066
rect 50410 87014 50422 87066
rect 50422 87014 50436 87066
rect 50460 87014 50474 87066
rect 50474 87014 50486 87066
rect 50486 87014 50516 87066
rect 50540 87014 50550 87066
rect 50550 87014 50596 87066
rect 50300 87012 50356 87014
rect 50380 87012 50436 87014
rect 50460 87012 50516 87014
rect 50540 87012 50596 87014
rect 50300 85978 50356 85980
rect 50380 85978 50436 85980
rect 50460 85978 50516 85980
rect 50540 85978 50596 85980
rect 50300 85926 50346 85978
rect 50346 85926 50356 85978
rect 50380 85926 50410 85978
rect 50410 85926 50422 85978
rect 50422 85926 50436 85978
rect 50460 85926 50474 85978
rect 50474 85926 50486 85978
rect 50486 85926 50516 85978
rect 50540 85926 50550 85978
rect 50550 85926 50596 85978
rect 50300 85924 50356 85926
rect 50380 85924 50436 85926
rect 50460 85924 50516 85926
rect 50540 85924 50596 85926
rect 50300 84890 50356 84892
rect 50380 84890 50436 84892
rect 50460 84890 50516 84892
rect 50540 84890 50596 84892
rect 50300 84838 50346 84890
rect 50346 84838 50356 84890
rect 50380 84838 50410 84890
rect 50410 84838 50422 84890
rect 50422 84838 50436 84890
rect 50460 84838 50474 84890
rect 50474 84838 50486 84890
rect 50486 84838 50516 84890
rect 50540 84838 50550 84890
rect 50550 84838 50596 84890
rect 50300 84836 50356 84838
rect 50380 84836 50436 84838
rect 50460 84836 50516 84838
rect 50540 84836 50596 84838
rect 50300 83802 50356 83804
rect 50380 83802 50436 83804
rect 50460 83802 50516 83804
rect 50540 83802 50596 83804
rect 50300 83750 50346 83802
rect 50346 83750 50356 83802
rect 50380 83750 50410 83802
rect 50410 83750 50422 83802
rect 50422 83750 50436 83802
rect 50460 83750 50474 83802
rect 50474 83750 50486 83802
rect 50486 83750 50516 83802
rect 50540 83750 50550 83802
rect 50550 83750 50596 83802
rect 50300 83748 50356 83750
rect 50380 83748 50436 83750
rect 50460 83748 50516 83750
rect 50540 83748 50596 83750
rect 50300 82714 50356 82716
rect 50380 82714 50436 82716
rect 50460 82714 50516 82716
rect 50540 82714 50596 82716
rect 50300 82662 50346 82714
rect 50346 82662 50356 82714
rect 50380 82662 50410 82714
rect 50410 82662 50422 82714
rect 50422 82662 50436 82714
rect 50460 82662 50474 82714
rect 50474 82662 50486 82714
rect 50486 82662 50516 82714
rect 50540 82662 50550 82714
rect 50550 82662 50596 82714
rect 50300 82660 50356 82662
rect 50380 82660 50436 82662
rect 50460 82660 50516 82662
rect 50540 82660 50596 82662
rect 50300 81626 50356 81628
rect 50380 81626 50436 81628
rect 50460 81626 50516 81628
rect 50540 81626 50596 81628
rect 50300 81574 50346 81626
rect 50346 81574 50356 81626
rect 50380 81574 50410 81626
rect 50410 81574 50422 81626
rect 50422 81574 50436 81626
rect 50460 81574 50474 81626
rect 50474 81574 50486 81626
rect 50486 81574 50516 81626
rect 50540 81574 50550 81626
rect 50550 81574 50596 81626
rect 50300 81572 50356 81574
rect 50380 81572 50436 81574
rect 50460 81572 50516 81574
rect 50540 81572 50596 81574
rect 50300 80538 50356 80540
rect 50380 80538 50436 80540
rect 50460 80538 50516 80540
rect 50540 80538 50596 80540
rect 50300 80486 50346 80538
rect 50346 80486 50356 80538
rect 50380 80486 50410 80538
rect 50410 80486 50422 80538
rect 50422 80486 50436 80538
rect 50460 80486 50474 80538
rect 50474 80486 50486 80538
rect 50486 80486 50516 80538
rect 50540 80486 50550 80538
rect 50550 80486 50596 80538
rect 50300 80484 50356 80486
rect 50380 80484 50436 80486
rect 50460 80484 50516 80486
rect 50540 80484 50596 80486
rect 50300 79450 50356 79452
rect 50380 79450 50436 79452
rect 50460 79450 50516 79452
rect 50540 79450 50596 79452
rect 50300 79398 50346 79450
rect 50346 79398 50356 79450
rect 50380 79398 50410 79450
rect 50410 79398 50422 79450
rect 50422 79398 50436 79450
rect 50460 79398 50474 79450
rect 50474 79398 50486 79450
rect 50486 79398 50516 79450
rect 50540 79398 50550 79450
rect 50550 79398 50596 79450
rect 50300 79396 50356 79398
rect 50380 79396 50436 79398
rect 50460 79396 50516 79398
rect 50540 79396 50596 79398
rect 50300 78362 50356 78364
rect 50380 78362 50436 78364
rect 50460 78362 50516 78364
rect 50540 78362 50596 78364
rect 50300 78310 50346 78362
rect 50346 78310 50356 78362
rect 50380 78310 50410 78362
rect 50410 78310 50422 78362
rect 50422 78310 50436 78362
rect 50460 78310 50474 78362
rect 50474 78310 50486 78362
rect 50486 78310 50516 78362
rect 50540 78310 50550 78362
rect 50550 78310 50596 78362
rect 50300 78308 50356 78310
rect 50380 78308 50436 78310
rect 50460 78308 50516 78310
rect 50540 78308 50596 78310
rect 50300 77274 50356 77276
rect 50380 77274 50436 77276
rect 50460 77274 50516 77276
rect 50540 77274 50596 77276
rect 50300 77222 50346 77274
rect 50346 77222 50356 77274
rect 50380 77222 50410 77274
rect 50410 77222 50422 77274
rect 50422 77222 50436 77274
rect 50460 77222 50474 77274
rect 50474 77222 50486 77274
rect 50486 77222 50516 77274
rect 50540 77222 50550 77274
rect 50550 77222 50596 77274
rect 50300 77220 50356 77222
rect 50380 77220 50436 77222
rect 50460 77220 50516 77222
rect 50540 77220 50596 77222
rect 50300 76186 50356 76188
rect 50380 76186 50436 76188
rect 50460 76186 50516 76188
rect 50540 76186 50596 76188
rect 50300 76134 50346 76186
rect 50346 76134 50356 76186
rect 50380 76134 50410 76186
rect 50410 76134 50422 76186
rect 50422 76134 50436 76186
rect 50460 76134 50474 76186
rect 50474 76134 50486 76186
rect 50486 76134 50516 76186
rect 50540 76134 50550 76186
rect 50550 76134 50596 76186
rect 50300 76132 50356 76134
rect 50380 76132 50436 76134
rect 50460 76132 50516 76134
rect 50540 76132 50596 76134
rect 50300 75098 50356 75100
rect 50380 75098 50436 75100
rect 50460 75098 50516 75100
rect 50540 75098 50596 75100
rect 50300 75046 50346 75098
rect 50346 75046 50356 75098
rect 50380 75046 50410 75098
rect 50410 75046 50422 75098
rect 50422 75046 50436 75098
rect 50460 75046 50474 75098
rect 50474 75046 50486 75098
rect 50486 75046 50516 75098
rect 50540 75046 50550 75098
rect 50550 75046 50596 75098
rect 50300 75044 50356 75046
rect 50380 75044 50436 75046
rect 50460 75044 50516 75046
rect 50540 75044 50596 75046
rect 50300 74010 50356 74012
rect 50380 74010 50436 74012
rect 50460 74010 50516 74012
rect 50540 74010 50596 74012
rect 50300 73958 50346 74010
rect 50346 73958 50356 74010
rect 50380 73958 50410 74010
rect 50410 73958 50422 74010
rect 50422 73958 50436 74010
rect 50460 73958 50474 74010
rect 50474 73958 50486 74010
rect 50486 73958 50516 74010
rect 50540 73958 50550 74010
rect 50550 73958 50596 74010
rect 50300 73956 50356 73958
rect 50380 73956 50436 73958
rect 50460 73956 50516 73958
rect 50540 73956 50596 73958
rect 50300 72922 50356 72924
rect 50380 72922 50436 72924
rect 50460 72922 50516 72924
rect 50540 72922 50596 72924
rect 50300 72870 50346 72922
rect 50346 72870 50356 72922
rect 50380 72870 50410 72922
rect 50410 72870 50422 72922
rect 50422 72870 50436 72922
rect 50460 72870 50474 72922
rect 50474 72870 50486 72922
rect 50486 72870 50516 72922
rect 50540 72870 50550 72922
rect 50550 72870 50596 72922
rect 50300 72868 50356 72870
rect 50380 72868 50436 72870
rect 50460 72868 50516 72870
rect 50540 72868 50596 72870
rect 50300 71834 50356 71836
rect 50380 71834 50436 71836
rect 50460 71834 50516 71836
rect 50540 71834 50596 71836
rect 50300 71782 50346 71834
rect 50346 71782 50356 71834
rect 50380 71782 50410 71834
rect 50410 71782 50422 71834
rect 50422 71782 50436 71834
rect 50460 71782 50474 71834
rect 50474 71782 50486 71834
rect 50486 71782 50516 71834
rect 50540 71782 50550 71834
rect 50550 71782 50596 71834
rect 50300 71780 50356 71782
rect 50380 71780 50436 71782
rect 50460 71780 50516 71782
rect 50540 71780 50596 71782
rect 50300 70746 50356 70748
rect 50380 70746 50436 70748
rect 50460 70746 50516 70748
rect 50540 70746 50596 70748
rect 50300 70694 50346 70746
rect 50346 70694 50356 70746
rect 50380 70694 50410 70746
rect 50410 70694 50422 70746
rect 50422 70694 50436 70746
rect 50460 70694 50474 70746
rect 50474 70694 50486 70746
rect 50486 70694 50516 70746
rect 50540 70694 50550 70746
rect 50550 70694 50596 70746
rect 50300 70692 50356 70694
rect 50380 70692 50436 70694
rect 50460 70692 50516 70694
rect 50540 70692 50596 70694
rect 50300 69658 50356 69660
rect 50380 69658 50436 69660
rect 50460 69658 50516 69660
rect 50540 69658 50596 69660
rect 50300 69606 50346 69658
rect 50346 69606 50356 69658
rect 50380 69606 50410 69658
rect 50410 69606 50422 69658
rect 50422 69606 50436 69658
rect 50460 69606 50474 69658
rect 50474 69606 50486 69658
rect 50486 69606 50516 69658
rect 50540 69606 50550 69658
rect 50550 69606 50596 69658
rect 50300 69604 50356 69606
rect 50380 69604 50436 69606
rect 50460 69604 50516 69606
rect 50540 69604 50596 69606
rect 50300 68570 50356 68572
rect 50380 68570 50436 68572
rect 50460 68570 50516 68572
rect 50540 68570 50596 68572
rect 50300 68518 50346 68570
rect 50346 68518 50356 68570
rect 50380 68518 50410 68570
rect 50410 68518 50422 68570
rect 50422 68518 50436 68570
rect 50460 68518 50474 68570
rect 50474 68518 50486 68570
rect 50486 68518 50516 68570
rect 50540 68518 50550 68570
rect 50550 68518 50596 68570
rect 50300 68516 50356 68518
rect 50380 68516 50436 68518
rect 50460 68516 50516 68518
rect 50540 68516 50596 68518
rect 50300 67482 50356 67484
rect 50380 67482 50436 67484
rect 50460 67482 50516 67484
rect 50540 67482 50596 67484
rect 50300 67430 50346 67482
rect 50346 67430 50356 67482
rect 50380 67430 50410 67482
rect 50410 67430 50422 67482
rect 50422 67430 50436 67482
rect 50460 67430 50474 67482
rect 50474 67430 50486 67482
rect 50486 67430 50516 67482
rect 50540 67430 50550 67482
rect 50550 67430 50596 67482
rect 50300 67428 50356 67430
rect 50380 67428 50436 67430
rect 50460 67428 50516 67430
rect 50540 67428 50596 67430
rect 50300 66394 50356 66396
rect 50380 66394 50436 66396
rect 50460 66394 50516 66396
rect 50540 66394 50596 66396
rect 50300 66342 50346 66394
rect 50346 66342 50356 66394
rect 50380 66342 50410 66394
rect 50410 66342 50422 66394
rect 50422 66342 50436 66394
rect 50460 66342 50474 66394
rect 50474 66342 50486 66394
rect 50486 66342 50516 66394
rect 50540 66342 50550 66394
rect 50550 66342 50596 66394
rect 50300 66340 50356 66342
rect 50380 66340 50436 66342
rect 50460 66340 50516 66342
rect 50540 66340 50596 66342
rect 50300 65306 50356 65308
rect 50380 65306 50436 65308
rect 50460 65306 50516 65308
rect 50540 65306 50596 65308
rect 50300 65254 50346 65306
rect 50346 65254 50356 65306
rect 50380 65254 50410 65306
rect 50410 65254 50422 65306
rect 50422 65254 50436 65306
rect 50460 65254 50474 65306
rect 50474 65254 50486 65306
rect 50486 65254 50516 65306
rect 50540 65254 50550 65306
rect 50550 65254 50596 65306
rect 50300 65252 50356 65254
rect 50380 65252 50436 65254
rect 50460 65252 50516 65254
rect 50540 65252 50596 65254
rect 50300 64218 50356 64220
rect 50380 64218 50436 64220
rect 50460 64218 50516 64220
rect 50540 64218 50596 64220
rect 50300 64166 50346 64218
rect 50346 64166 50356 64218
rect 50380 64166 50410 64218
rect 50410 64166 50422 64218
rect 50422 64166 50436 64218
rect 50460 64166 50474 64218
rect 50474 64166 50486 64218
rect 50486 64166 50516 64218
rect 50540 64166 50550 64218
rect 50550 64166 50596 64218
rect 50300 64164 50356 64166
rect 50380 64164 50436 64166
rect 50460 64164 50516 64166
rect 50540 64164 50596 64166
rect 50300 63130 50356 63132
rect 50380 63130 50436 63132
rect 50460 63130 50516 63132
rect 50540 63130 50596 63132
rect 50300 63078 50346 63130
rect 50346 63078 50356 63130
rect 50380 63078 50410 63130
rect 50410 63078 50422 63130
rect 50422 63078 50436 63130
rect 50460 63078 50474 63130
rect 50474 63078 50486 63130
rect 50486 63078 50516 63130
rect 50540 63078 50550 63130
rect 50550 63078 50596 63130
rect 50300 63076 50356 63078
rect 50380 63076 50436 63078
rect 50460 63076 50516 63078
rect 50540 63076 50596 63078
rect 50300 62042 50356 62044
rect 50380 62042 50436 62044
rect 50460 62042 50516 62044
rect 50540 62042 50596 62044
rect 50300 61990 50346 62042
rect 50346 61990 50356 62042
rect 50380 61990 50410 62042
rect 50410 61990 50422 62042
rect 50422 61990 50436 62042
rect 50460 61990 50474 62042
rect 50474 61990 50486 62042
rect 50486 61990 50516 62042
rect 50540 61990 50550 62042
rect 50550 61990 50596 62042
rect 50300 61988 50356 61990
rect 50380 61988 50436 61990
rect 50460 61988 50516 61990
rect 50540 61988 50596 61990
rect 50300 60954 50356 60956
rect 50380 60954 50436 60956
rect 50460 60954 50516 60956
rect 50540 60954 50596 60956
rect 50300 60902 50346 60954
rect 50346 60902 50356 60954
rect 50380 60902 50410 60954
rect 50410 60902 50422 60954
rect 50422 60902 50436 60954
rect 50460 60902 50474 60954
rect 50474 60902 50486 60954
rect 50486 60902 50516 60954
rect 50540 60902 50550 60954
rect 50550 60902 50596 60954
rect 50300 60900 50356 60902
rect 50380 60900 50436 60902
rect 50460 60900 50516 60902
rect 50540 60900 50596 60902
rect 50300 59866 50356 59868
rect 50380 59866 50436 59868
rect 50460 59866 50516 59868
rect 50540 59866 50596 59868
rect 50300 59814 50346 59866
rect 50346 59814 50356 59866
rect 50380 59814 50410 59866
rect 50410 59814 50422 59866
rect 50422 59814 50436 59866
rect 50460 59814 50474 59866
rect 50474 59814 50486 59866
rect 50486 59814 50516 59866
rect 50540 59814 50550 59866
rect 50550 59814 50596 59866
rect 50300 59812 50356 59814
rect 50380 59812 50436 59814
rect 50460 59812 50516 59814
rect 50540 59812 50596 59814
rect 50300 58778 50356 58780
rect 50380 58778 50436 58780
rect 50460 58778 50516 58780
rect 50540 58778 50596 58780
rect 50300 58726 50346 58778
rect 50346 58726 50356 58778
rect 50380 58726 50410 58778
rect 50410 58726 50422 58778
rect 50422 58726 50436 58778
rect 50460 58726 50474 58778
rect 50474 58726 50486 58778
rect 50486 58726 50516 58778
rect 50540 58726 50550 58778
rect 50550 58726 50596 58778
rect 50300 58724 50356 58726
rect 50380 58724 50436 58726
rect 50460 58724 50516 58726
rect 50540 58724 50596 58726
rect 50300 57690 50356 57692
rect 50380 57690 50436 57692
rect 50460 57690 50516 57692
rect 50540 57690 50596 57692
rect 50300 57638 50346 57690
rect 50346 57638 50356 57690
rect 50380 57638 50410 57690
rect 50410 57638 50422 57690
rect 50422 57638 50436 57690
rect 50460 57638 50474 57690
rect 50474 57638 50486 57690
rect 50486 57638 50516 57690
rect 50540 57638 50550 57690
rect 50550 57638 50596 57690
rect 50300 57636 50356 57638
rect 50380 57636 50436 57638
rect 50460 57636 50516 57638
rect 50540 57636 50596 57638
rect 50300 56602 50356 56604
rect 50380 56602 50436 56604
rect 50460 56602 50516 56604
rect 50540 56602 50596 56604
rect 50300 56550 50346 56602
rect 50346 56550 50356 56602
rect 50380 56550 50410 56602
rect 50410 56550 50422 56602
rect 50422 56550 50436 56602
rect 50460 56550 50474 56602
rect 50474 56550 50486 56602
rect 50486 56550 50516 56602
rect 50540 56550 50550 56602
rect 50550 56550 50596 56602
rect 50300 56548 50356 56550
rect 50380 56548 50436 56550
rect 50460 56548 50516 56550
rect 50540 56548 50596 56550
rect 50300 55514 50356 55516
rect 50380 55514 50436 55516
rect 50460 55514 50516 55516
rect 50540 55514 50596 55516
rect 50300 55462 50346 55514
rect 50346 55462 50356 55514
rect 50380 55462 50410 55514
rect 50410 55462 50422 55514
rect 50422 55462 50436 55514
rect 50460 55462 50474 55514
rect 50474 55462 50486 55514
rect 50486 55462 50516 55514
rect 50540 55462 50550 55514
rect 50550 55462 50596 55514
rect 50300 55460 50356 55462
rect 50380 55460 50436 55462
rect 50460 55460 50516 55462
rect 50540 55460 50596 55462
rect 50300 54426 50356 54428
rect 50380 54426 50436 54428
rect 50460 54426 50516 54428
rect 50540 54426 50596 54428
rect 50300 54374 50346 54426
rect 50346 54374 50356 54426
rect 50380 54374 50410 54426
rect 50410 54374 50422 54426
rect 50422 54374 50436 54426
rect 50460 54374 50474 54426
rect 50474 54374 50486 54426
rect 50486 54374 50516 54426
rect 50540 54374 50550 54426
rect 50550 54374 50596 54426
rect 50300 54372 50356 54374
rect 50380 54372 50436 54374
rect 50460 54372 50516 54374
rect 50540 54372 50596 54374
rect 50300 53338 50356 53340
rect 50380 53338 50436 53340
rect 50460 53338 50516 53340
rect 50540 53338 50596 53340
rect 50300 53286 50346 53338
rect 50346 53286 50356 53338
rect 50380 53286 50410 53338
rect 50410 53286 50422 53338
rect 50422 53286 50436 53338
rect 50460 53286 50474 53338
rect 50474 53286 50486 53338
rect 50486 53286 50516 53338
rect 50540 53286 50550 53338
rect 50550 53286 50596 53338
rect 50300 53284 50356 53286
rect 50380 53284 50436 53286
rect 50460 53284 50516 53286
rect 50540 53284 50596 53286
rect 50300 52250 50356 52252
rect 50380 52250 50436 52252
rect 50460 52250 50516 52252
rect 50540 52250 50596 52252
rect 50300 52198 50346 52250
rect 50346 52198 50356 52250
rect 50380 52198 50410 52250
rect 50410 52198 50422 52250
rect 50422 52198 50436 52250
rect 50460 52198 50474 52250
rect 50474 52198 50486 52250
rect 50486 52198 50516 52250
rect 50540 52198 50550 52250
rect 50550 52198 50596 52250
rect 50300 52196 50356 52198
rect 50380 52196 50436 52198
rect 50460 52196 50516 52198
rect 50540 52196 50596 52198
rect 50300 51162 50356 51164
rect 50380 51162 50436 51164
rect 50460 51162 50516 51164
rect 50540 51162 50596 51164
rect 50300 51110 50346 51162
rect 50346 51110 50356 51162
rect 50380 51110 50410 51162
rect 50410 51110 50422 51162
rect 50422 51110 50436 51162
rect 50460 51110 50474 51162
rect 50474 51110 50486 51162
rect 50486 51110 50516 51162
rect 50540 51110 50550 51162
rect 50550 51110 50596 51162
rect 50300 51108 50356 51110
rect 50380 51108 50436 51110
rect 50460 51108 50516 51110
rect 50540 51108 50596 51110
rect 50300 50074 50356 50076
rect 50380 50074 50436 50076
rect 50460 50074 50516 50076
rect 50540 50074 50596 50076
rect 50300 50022 50346 50074
rect 50346 50022 50356 50074
rect 50380 50022 50410 50074
rect 50410 50022 50422 50074
rect 50422 50022 50436 50074
rect 50460 50022 50474 50074
rect 50474 50022 50486 50074
rect 50486 50022 50516 50074
rect 50540 50022 50550 50074
rect 50550 50022 50596 50074
rect 50300 50020 50356 50022
rect 50380 50020 50436 50022
rect 50460 50020 50516 50022
rect 50540 50020 50596 50022
rect 50300 48986 50356 48988
rect 50380 48986 50436 48988
rect 50460 48986 50516 48988
rect 50540 48986 50596 48988
rect 50300 48934 50346 48986
rect 50346 48934 50356 48986
rect 50380 48934 50410 48986
rect 50410 48934 50422 48986
rect 50422 48934 50436 48986
rect 50460 48934 50474 48986
rect 50474 48934 50486 48986
rect 50486 48934 50516 48986
rect 50540 48934 50550 48986
rect 50550 48934 50596 48986
rect 50300 48932 50356 48934
rect 50380 48932 50436 48934
rect 50460 48932 50516 48934
rect 50540 48932 50596 48934
rect 50300 47898 50356 47900
rect 50380 47898 50436 47900
rect 50460 47898 50516 47900
rect 50540 47898 50596 47900
rect 50300 47846 50346 47898
rect 50346 47846 50356 47898
rect 50380 47846 50410 47898
rect 50410 47846 50422 47898
rect 50422 47846 50436 47898
rect 50460 47846 50474 47898
rect 50474 47846 50486 47898
rect 50486 47846 50516 47898
rect 50540 47846 50550 47898
rect 50550 47846 50596 47898
rect 50300 47844 50356 47846
rect 50380 47844 50436 47846
rect 50460 47844 50516 47846
rect 50540 47844 50596 47846
rect 50300 46810 50356 46812
rect 50380 46810 50436 46812
rect 50460 46810 50516 46812
rect 50540 46810 50596 46812
rect 50300 46758 50346 46810
rect 50346 46758 50356 46810
rect 50380 46758 50410 46810
rect 50410 46758 50422 46810
rect 50422 46758 50436 46810
rect 50460 46758 50474 46810
rect 50474 46758 50486 46810
rect 50486 46758 50516 46810
rect 50540 46758 50550 46810
rect 50550 46758 50596 46810
rect 50300 46756 50356 46758
rect 50380 46756 50436 46758
rect 50460 46756 50516 46758
rect 50540 46756 50596 46758
rect 50300 45722 50356 45724
rect 50380 45722 50436 45724
rect 50460 45722 50516 45724
rect 50540 45722 50596 45724
rect 50300 45670 50346 45722
rect 50346 45670 50356 45722
rect 50380 45670 50410 45722
rect 50410 45670 50422 45722
rect 50422 45670 50436 45722
rect 50460 45670 50474 45722
rect 50474 45670 50486 45722
rect 50486 45670 50516 45722
rect 50540 45670 50550 45722
rect 50550 45670 50596 45722
rect 50300 45668 50356 45670
rect 50380 45668 50436 45670
rect 50460 45668 50516 45670
rect 50540 45668 50596 45670
rect 50300 44634 50356 44636
rect 50380 44634 50436 44636
rect 50460 44634 50516 44636
rect 50540 44634 50596 44636
rect 50300 44582 50346 44634
rect 50346 44582 50356 44634
rect 50380 44582 50410 44634
rect 50410 44582 50422 44634
rect 50422 44582 50436 44634
rect 50460 44582 50474 44634
rect 50474 44582 50486 44634
rect 50486 44582 50516 44634
rect 50540 44582 50550 44634
rect 50550 44582 50596 44634
rect 50300 44580 50356 44582
rect 50380 44580 50436 44582
rect 50460 44580 50516 44582
rect 50540 44580 50596 44582
rect 50300 43546 50356 43548
rect 50380 43546 50436 43548
rect 50460 43546 50516 43548
rect 50540 43546 50596 43548
rect 50300 43494 50346 43546
rect 50346 43494 50356 43546
rect 50380 43494 50410 43546
rect 50410 43494 50422 43546
rect 50422 43494 50436 43546
rect 50460 43494 50474 43546
rect 50474 43494 50486 43546
rect 50486 43494 50516 43546
rect 50540 43494 50550 43546
rect 50550 43494 50596 43546
rect 50300 43492 50356 43494
rect 50380 43492 50436 43494
rect 50460 43492 50516 43494
rect 50540 43492 50596 43494
rect 50300 42458 50356 42460
rect 50380 42458 50436 42460
rect 50460 42458 50516 42460
rect 50540 42458 50596 42460
rect 50300 42406 50346 42458
rect 50346 42406 50356 42458
rect 50380 42406 50410 42458
rect 50410 42406 50422 42458
rect 50422 42406 50436 42458
rect 50460 42406 50474 42458
rect 50474 42406 50486 42458
rect 50486 42406 50516 42458
rect 50540 42406 50550 42458
rect 50550 42406 50596 42458
rect 50300 42404 50356 42406
rect 50380 42404 50436 42406
rect 50460 42404 50516 42406
rect 50540 42404 50596 42406
rect 50300 41370 50356 41372
rect 50380 41370 50436 41372
rect 50460 41370 50516 41372
rect 50540 41370 50596 41372
rect 50300 41318 50346 41370
rect 50346 41318 50356 41370
rect 50380 41318 50410 41370
rect 50410 41318 50422 41370
rect 50422 41318 50436 41370
rect 50460 41318 50474 41370
rect 50474 41318 50486 41370
rect 50486 41318 50516 41370
rect 50540 41318 50550 41370
rect 50550 41318 50596 41370
rect 50300 41316 50356 41318
rect 50380 41316 50436 41318
rect 50460 41316 50516 41318
rect 50540 41316 50596 41318
rect 50300 40282 50356 40284
rect 50380 40282 50436 40284
rect 50460 40282 50516 40284
rect 50540 40282 50596 40284
rect 50300 40230 50346 40282
rect 50346 40230 50356 40282
rect 50380 40230 50410 40282
rect 50410 40230 50422 40282
rect 50422 40230 50436 40282
rect 50460 40230 50474 40282
rect 50474 40230 50486 40282
rect 50486 40230 50516 40282
rect 50540 40230 50550 40282
rect 50550 40230 50596 40282
rect 50300 40228 50356 40230
rect 50380 40228 50436 40230
rect 50460 40228 50516 40230
rect 50540 40228 50596 40230
rect 50300 39194 50356 39196
rect 50380 39194 50436 39196
rect 50460 39194 50516 39196
rect 50540 39194 50596 39196
rect 50300 39142 50346 39194
rect 50346 39142 50356 39194
rect 50380 39142 50410 39194
rect 50410 39142 50422 39194
rect 50422 39142 50436 39194
rect 50460 39142 50474 39194
rect 50474 39142 50486 39194
rect 50486 39142 50516 39194
rect 50540 39142 50550 39194
rect 50550 39142 50596 39194
rect 50300 39140 50356 39142
rect 50380 39140 50436 39142
rect 50460 39140 50516 39142
rect 50540 39140 50596 39142
rect 50300 38106 50356 38108
rect 50380 38106 50436 38108
rect 50460 38106 50516 38108
rect 50540 38106 50596 38108
rect 50300 38054 50346 38106
rect 50346 38054 50356 38106
rect 50380 38054 50410 38106
rect 50410 38054 50422 38106
rect 50422 38054 50436 38106
rect 50460 38054 50474 38106
rect 50474 38054 50486 38106
rect 50486 38054 50516 38106
rect 50540 38054 50550 38106
rect 50550 38054 50596 38106
rect 50300 38052 50356 38054
rect 50380 38052 50436 38054
rect 50460 38052 50516 38054
rect 50540 38052 50596 38054
rect 50300 37018 50356 37020
rect 50380 37018 50436 37020
rect 50460 37018 50516 37020
rect 50540 37018 50596 37020
rect 50300 36966 50346 37018
rect 50346 36966 50356 37018
rect 50380 36966 50410 37018
rect 50410 36966 50422 37018
rect 50422 36966 50436 37018
rect 50460 36966 50474 37018
rect 50474 36966 50486 37018
rect 50486 36966 50516 37018
rect 50540 36966 50550 37018
rect 50550 36966 50596 37018
rect 50300 36964 50356 36966
rect 50380 36964 50436 36966
rect 50460 36964 50516 36966
rect 50540 36964 50596 36966
rect 50300 35930 50356 35932
rect 50380 35930 50436 35932
rect 50460 35930 50516 35932
rect 50540 35930 50596 35932
rect 50300 35878 50346 35930
rect 50346 35878 50356 35930
rect 50380 35878 50410 35930
rect 50410 35878 50422 35930
rect 50422 35878 50436 35930
rect 50460 35878 50474 35930
rect 50474 35878 50486 35930
rect 50486 35878 50516 35930
rect 50540 35878 50550 35930
rect 50550 35878 50596 35930
rect 50300 35876 50356 35878
rect 50380 35876 50436 35878
rect 50460 35876 50516 35878
rect 50540 35876 50596 35878
rect 50300 34842 50356 34844
rect 50380 34842 50436 34844
rect 50460 34842 50516 34844
rect 50540 34842 50596 34844
rect 50300 34790 50346 34842
rect 50346 34790 50356 34842
rect 50380 34790 50410 34842
rect 50410 34790 50422 34842
rect 50422 34790 50436 34842
rect 50460 34790 50474 34842
rect 50474 34790 50486 34842
rect 50486 34790 50516 34842
rect 50540 34790 50550 34842
rect 50550 34790 50596 34842
rect 50300 34788 50356 34790
rect 50380 34788 50436 34790
rect 50460 34788 50516 34790
rect 50540 34788 50596 34790
rect 50300 33754 50356 33756
rect 50380 33754 50436 33756
rect 50460 33754 50516 33756
rect 50540 33754 50596 33756
rect 50300 33702 50346 33754
rect 50346 33702 50356 33754
rect 50380 33702 50410 33754
rect 50410 33702 50422 33754
rect 50422 33702 50436 33754
rect 50460 33702 50474 33754
rect 50474 33702 50486 33754
rect 50486 33702 50516 33754
rect 50540 33702 50550 33754
rect 50550 33702 50596 33754
rect 50300 33700 50356 33702
rect 50380 33700 50436 33702
rect 50460 33700 50516 33702
rect 50540 33700 50596 33702
rect 50300 32666 50356 32668
rect 50380 32666 50436 32668
rect 50460 32666 50516 32668
rect 50540 32666 50596 32668
rect 50300 32614 50346 32666
rect 50346 32614 50356 32666
rect 50380 32614 50410 32666
rect 50410 32614 50422 32666
rect 50422 32614 50436 32666
rect 50460 32614 50474 32666
rect 50474 32614 50486 32666
rect 50486 32614 50516 32666
rect 50540 32614 50550 32666
rect 50550 32614 50596 32666
rect 50300 32612 50356 32614
rect 50380 32612 50436 32614
rect 50460 32612 50516 32614
rect 50540 32612 50596 32614
rect 50300 31578 50356 31580
rect 50380 31578 50436 31580
rect 50460 31578 50516 31580
rect 50540 31578 50596 31580
rect 50300 31526 50346 31578
rect 50346 31526 50356 31578
rect 50380 31526 50410 31578
rect 50410 31526 50422 31578
rect 50422 31526 50436 31578
rect 50460 31526 50474 31578
rect 50474 31526 50486 31578
rect 50486 31526 50516 31578
rect 50540 31526 50550 31578
rect 50550 31526 50596 31578
rect 50300 31524 50356 31526
rect 50380 31524 50436 31526
rect 50460 31524 50516 31526
rect 50540 31524 50596 31526
rect 50300 30490 50356 30492
rect 50380 30490 50436 30492
rect 50460 30490 50516 30492
rect 50540 30490 50596 30492
rect 50300 30438 50346 30490
rect 50346 30438 50356 30490
rect 50380 30438 50410 30490
rect 50410 30438 50422 30490
rect 50422 30438 50436 30490
rect 50460 30438 50474 30490
rect 50474 30438 50486 30490
rect 50486 30438 50516 30490
rect 50540 30438 50550 30490
rect 50550 30438 50596 30490
rect 50300 30436 50356 30438
rect 50380 30436 50436 30438
rect 50460 30436 50516 30438
rect 50540 30436 50596 30438
rect 50300 29402 50356 29404
rect 50380 29402 50436 29404
rect 50460 29402 50516 29404
rect 50540 29402 50596 29404
rect 50300 29350 50346 29402
rect 50346 29350 50356 29402
rect 50380 29350 50410 29402
rect 50410 29350 50422 29402
rect 50422 29350 50436 29402
rect 50460 29350 50474 29402
rect 50474 29350 50486 29402
rect 50486 29350 50516 29402
rect 50540 29350 50550 29402
rect 50550 29350 50596 29402
rect 50300 29348 50356 29350
rect 50380 29348 50436 29350
rect 50460 29348 50516 29350
rect 50540 29348 50596 29350
rect 50300 28314 50356 28316
rect 50380 28314 50436 28316
rect 50460 28314 50516 28316
rect 50540 28314 50596 28316
rect 50300 28262 50346 28314
rect 50346 28262 50356 28314
rect 50380 28262 50410 28314
rect 50410 28262 50422 28314
rect 50422 28262 50436 28314
rect 50460 28262 50474 28314
rect 50474 28262 50486 28314
rect 50486 28262 50516 28314
rect 50540 28262 50550 28314
rect 50550 28262 50596 28314
rect 50300 28260 50356 28262
rect 50380 28260 50436 28262
rect 50460 28260 50516 28262
rect 50540 28260 50596 28262
rect 50300 27226 50356 27228
rect 50380 27226 50436 27228
rect 50460 27226 50516 27228
rect 50540 27226 50596 27228
rect 50300 27174 50346 27226
rect 50346 27174 50356 27226
rect 50380 27174 50410 27226
rect 50410 27174 50422 27226
rect 50422 27174 50436 27226
rect 50460 27174 50474 27226
rect 50474 27174 50486 27226
rect 50486 27174 50516 27226
rect 50540 27174 50550 27226
rect 50550 27174 50596 27226
rect 50300 27172 50356 27174
rect 50380 27172 50436 27174
rect 50460 27172 50516 27174
rect 50540 27172 50596 27174
rect 50300 26138 50356 26140
rect 50380 26138 50436 26140
rect 50460 26138 50516 26140
rect 50540 26138 50596 26140
rect 50300 26086 50346 26138
rect 50346 26086 50356 26138
rect 50380 26086 50410 26138
rect 50410 26086 50422 26138
rect 50422 26086 50436 26138
rect 50460 26086 50474 26138
rect 50474 26086 50486 26138
rect 50486 26086 50516 26138
rect 50540 26086 50550 26138
rect 50550 26086 50596 26138
rect 50300 26084 50356 26086
rect 50380 26084 50436 26086
rect 50460 26084 50516 26086
rect 50540 26084 50596 26086
rect 50300 25050 50356 25052
rect 50380 25050 50436 25052
rect 50460 25050 50516 25052
rect 50540 25050 50596 25052
rect 50300 24998 50346 25050
rect 50346 24998 50356 25050
rect 50380 24998 50410 25050
rect 50410 24998 50422 25050
rect 50422 24998 50436 25050
rect 50460 24998 50474 25050
rect 50474 24998 50486 25050
rect 50486 24998 50516 25050
rect 50540 24998 50550 25050
rect 50550 24998 50596 25050
rect 50300 24996 50356 24998
rect 50380 24996 50436 24998
rect 50460 24996 50516 24998
rect 50540 24996 50596 24998
rect 50300 23962 50356 23964
rect 50380 23962 50436 23964
rect 50460 23962 50516 23964
rect 50540 23962 50596 23964
rect 50300 23910 50346 23962
rect 50346 23910 50356 23962
rect 50380 23910 50410 23962
rect 50410 23910 50422 23962
rect 50422 23910 50436 23962
rect 50460 23910 50474 23962
rect 50474 23910 50486 23962
rect 50486 23910 50516 23962
rect 50540 23910 50550 23962
rect 50550 23910 50596 23962
rect 50300 23908 50356 23910
rect 50380 23908 50436 23910
rect 50460 23908 50516 23910
rect 50540 23908 50596 23910
rect 50300 22874 50356 22876
rect 50380 22874 50436 22876
rect 50460 22874 50516 22876
rect 50540 22874 50596 22876
rect 50300 22822 50346 22874
rect 50346 22822 50356 22874
rect 50380 22822 50410 22874
rect 50410 22822 50422 22874
rect 50422 22822 50436 22874
rect 50460 22822 50474 22874
rect 50474 22822 50486 22874
rect 50486 22822 50516 22874
rect 50540 22822 50550 22874
rect 50550 22822 50596 22874
rect 50300 22820 50356 22822
rect 50380 22820 50436 22822
rect 50460 22820 50516 22822
rect 50540 22820 50596 22822
rect 50300 21786 50356 21788
rect 50380 21786 50436 21788
rect 50460 21786 50516 21788
rect 50540 21786 50596 21788
rect 50300 21734 50346 21786
rect 50346 21734 50356 21786
rect 50380 21734 50410 21786
rect 50410 21734 50422 21786
rect 50422 21734 50436 21786
rect 50460 21734 50474 21786
rect 50474 21734 50486 21786
rect 50486 21734 50516 21786
rect 50540 21734 50550 21786
rect 50550 21734 50596 21786
rect 50300 21732 50356 21734
rect 50380 21732 50436 21734
rect 50460 21732 50516 21734
rect 50540 21732 50596 21734
rect 50300 20698 50356 20700
rect 50380 20698 50436 20700
rect 50460 20698 50516 20700
rect 50540 20698 50596 20700
rect 50300 20646 50346 20698
rect 50346 20646 50356 20698
rect 50380 20646 50410 20698
rect 50410 20646 50422 20698
rect 50422 20646 50436 20698
rect 50460 20646 50474 20698
rect 50474 20646 50486 20698
rect 50486 20646 50516 20698
rect 50540 20646 50550 20698
rect 50550 20646 50596 20698
rect 50300 20644 50356 20646
rect 50380 20644 50436 20646
rect 50460 20644 50516 20646
rect 50540 20644 50596 20646
rect 50300 19610 50356 19612
rect 50380 19610 50436 19612
rect 50460 19610 50516 19612
rect 50540 19610 50596 19612
rect 50300 19558 50346 19610
rect 50346 19558 50356 19610
rect 50380 19558 50410 19610
rect 50410 19558 50422 19610
rect 50422 19558 50436 19610
rect 50460 19558 50474 19610
rect 50474 19558 50486 19610
rect 50486 19558 50516 19610
rect 50540 19558 50550 19610
rect 50550 19558 50596 19610
rect 50300 19556 50356 19558
rect 50380 19556 50436 19558
rect 50460 19556 50516 19558
rect 50540 19556 50596 19558
rect 50300 18522 50356 18524
rect 50380 18522 50436 18524
rect 50460 18522 50516 18524
rect 50540 18522 50596 18524
rect 50300 18470 50346 18522
rect 50346 18470 50356 18522
rect 50380 18470 50410 18522
rect 50410 18470 50422 18522
rect 50422 18470 50436 18522
rect 50460 18470 50474 18522
rect 50474 18470 50486 18522
rect 50486 18470 50516 18522
rect 50540 18470 50550 18522
rect 50550 18470 50596 18522
rect 50300 18468 50356 18470
rect 50380 18468 50436 18470
rect 50460 18468 50516 18470
rect 50540 18468 50596 18470
rect 50300 17434 50356 17436
rect 50380 17434 50436 17436
rect 50460 17434 50516 17436
rect 50540 17434 50596 17436
rect 50300 17382 50346 17434
rect 50346 17382 50356 17434
rect 50380 17382 50410 17434
rect 50410 17382 50422 17434
rect 50422 17382 50436 17434
rect 50460 17382 50474 17434
rect 50474 17382 50486 17434
rect 50486 17382 50516 17434
rect 50540 17382 50550 17434
rect 50550 17382 50596 17434
rect 50300 17380 50356 17382
rect 50380 17380 50436 17382
rect 50460 17380 50516 17382
rect 50540 17380 50596 17382
rect 77206 118360 77262 118416
rect 65660 116986 65716 116988
rect 65740 116986 65796 116988
rect 65820 116986 65876 116988
rect 65900 116986 65956 116988
rect 65660 116934 65706 116986
rect 65706 116934 65716 116986
rect 65740 116934 65770 116986
rect 65770 116934 65782 116986
rect 65782 116934 65796 116986
rect 65820 116934 65834 116986
rect 65834 116934 65846 116986
rect 65846 116934 65876 116986
rect 65900 116934 65910 116986
rect 65910 116934 65956 116986
rect 65660 116932 65716 116934
rect 65740 116932 65796 116934
rect 65820 116932 65876 116934
rect 65900 116932 65956 116934
rect 65660 115898 65716 115900
rect 65740 115898 65796 115900
rect 65820 115898 65876 115900
rect 65900 115898 65956 115900
rect 65660 115846 65706 115898
rect 65706 115846 65716 115898
rect 65740 115846 65770 115898
rect 65770 115846 65782 115898
rect 65782 115846 65796 115898
rect 65820 115846 65834 115898
rect 65834 115846 65846 115898
rect 65846 115846 65876 115898
rect 65900 115846 65910 115898
rect 65910 115846 65956 115898
rect 65660 115844 65716 115846
rect 65740 115844 65796 115846
rect 65820 115844 65876 115846
rect 65900 115844 65956 115846
rect 65660 114810 65716 114812
rect 65740 114810 65796 114812
rect 65820 114810 65876 114812
rect 65900 114810 65956 114812
rect 65660 114758 65706 114810
rect 65706 114758 65716 114810
rect 65740 114758 65770 114810
rect 65770 114758 65782 114810
rect 65782 114758 65796 114810
rect 65820 114758 65834 114810
rect 65834 114758 65846 114810
rect 65846 114758 65876 114810
rect 65900 114758 65910 114810
rect 65910 114758 65956 114810
rect 65660 114756 65716 114758
rect 65740 114756 65796 114758
rect 65820 114756 65876 114758
rect 65900 114756 65956 114758
rect 65660 113722 65716 113724
rect 65740 113722 65796 113724
rect 65820 113722 65876 113724
rect 65900 113722 65956 113724
rect 65660 113670 65706 113722
rect 65706 113670 65716 113722
rect 65740 113670 65770 113722
rect 65770 113670 65782 113722
rect 65782 113670 65796 113722
rect 65820 113670 65834 113722
rect 65834 113670 65846 113722
rect 65846 113670 65876 113722
rect 65900 113670 65910 113722
rect 65910 113670 65956 113722
rect 65660 113668 65716 113670
rect 65740 113668 65796 113670
rect 65820 113668 65876 113670
rect 65900 113668 65956 113670
rect 65660 112634 65716 112636
rect 65740 112634 65796 112636
rect 65820 112634 65876 112636
rect 65900 112634 65956 112636
rect 65660 112582 65706 112634
rect 65706 112582 65716 112634
rect 65740 112582 65770 112634
rect 65770 112582 65782 112634
rect 65782 112582 65796 112634
rect 65820 112582 65834 112634
rect 65834 112582 65846 112634
rect 65846 112582 65876 112634
rect 65900 112582 65910 112634
rect 65910 112582 65956 112634
rect 65660 112580 65716 112582
rect 65740 112580 65796 112582
rect 65820 112580 65876 112582
rect 65900 112580 65956 112582
rect 65660 111546 65716 111548
rect 65740 111546 65796 111548
rect 65820 111546 65876 111548
rect 65900 111546 65956 111548
rect 65660 111494 65706 111546
rect 65706 111494 65716 111546
rect 65740 111494 65770 111546
rect 65770 111494 65782 111546
rect 65782 111494 65796 111546
rect 65820 111494 65834 111546
rect 65834 111494 65846 111546
rect 65846 111494 65876 111546
rect 65900 111494 65910 111546
rect 65910 111494 65956 111546
rect 65660 111492 65716 111494
rect 65740 111492 65796 111494
rect 65820 111492 65876 111494
rect 65900 111492 65956 111494
rect 65660 110458 65716 110460
rect 65740 110458 65796 110460
rect 65820 110458 65876 110460
rect 65900 110458 65956 110460
rect 65660 110406 65706 110458
rect 65706 110406 65716 110458
rect 65740 110406 65770 110458
rect 65770 110406 65782 110458
rect 65782 110406 65796 110458
rect 65820 110406 65834 110458
rect 65834 110406 65846 110458
rect 65846 110406 65876 110458
rect 65900 110406 65910 110458
rect 65910 110406 65956 110458
rect 65660 110404 65716 110406
rect 65740 110404 65796 110406
rect 65820 110404 65876 110406
rect 65900 110404 65956 110406
rect 65660 109370 65716 109372
rect 65740 109370 65796 109372
rect 65820 109370 65876 109372
rect 65900 109370 65956 109372
rect 65660 109318 65706 109370
rect 65706 109318 65716 109370
rect 65740 109318 65770 109370
rect 65770 109318 65782 109370
rect 65782 109318 65796 109370
rect 65820 109318 65834 109370
rect 65834 109318 65846 109370
rect 65846 109318 65876 109370
rect 65900 109318 65910 109370
rect 65910 109318 65956 109370
rect 65660 109316 65716 109318
rect 65740 109316 65796 109318
rect 65820 109316 65876 109318
rect 65900 109316 65956 109318
rect 65660 108282 65716 108284
rect 65740 108282 65796 108284
rect 65820 108282 65876 108284
rect 65900 108282 65956 108284
rect 65660 108230 65706 108282
rect 65706 108230 65716 108282
rect 65740 108230 65770 108282
rect 65770 108230 65782 108282
rect 65782 108230 65796 108282
rect 65820 108230 65834 108282
rect 65834 108230 65846 108282
rect 65846 108230 65876 108282
rect 65900 108230 65910 108282
rect 65910 108230 65956 108282
rect 65660 108228 65716 108230
rect 65740 108228 65796 108230
rect 65820 108228 65876 108230
rect 65900 108228 65956 108230
rect 65660 107194 65716 107196
rect 65740 107194 65796 107196
rect 65820 107194 65876 107196
rect 65900 107194 65956 107196
rect 65660 107142 65706 107194
rect 65706 107142 65716 107194
rect 65740 107142 65770 107194
rect 65770 107142 65782 107194
rect 65782 107142 65796 107194
rect 65820 107142 65834 107194
rect 65834 107142 65846 107194
rect 65846 107142 65876 107194
rect 65900 107142 65910 107194
rect 65910 107142 65956 107194
rect 65660 107140 65716 107142
rect 65740 107140 65796 107142
rect 65820 107140 65876 107142
rect 65900 107140 65956 107142
rect 65660 106106 65716 106108
rect 65740 106106 65796 106108
rect 65820 106106 65876 106108
rect 65900 106106 65956 106108
rect 65660 106054 65706 106106
rect 65706 106054 65716 106106
rect 65740 106054 65770 106106
rect 65770 106054 65782 106106
rect 65782 106054 65796 106106
rect 65820 106054 65834 106106
rect 65834 106054 65846 106106
rect 65846 106054 65876 106106
rect 65900 106054 65910 106106
rect 65910 106054 65956 106106
rect 65660 106052 65716 106054
rect 65740 106052 65796 106054
rect 65820 106052 65876 106054
rect 65900 106052 65956 106054
rect 65660 105018 65716 105020
rect 65740 105018 65796 105020
rect 65820 105018 65876 105020
rect 65900 105018 65956 105020
rect 65660 104966 65706 105018
rect 65706 104966 65716 105018
rect 65740 104966 65770 105018
rect 65770 104966 65782 105018
rect 65782 104966 65796 105018
rect 65820 104966 65834 105018
rect 65834 104966 65846 105018
rect 65846 104966 65876 105018
rect 65900 104966 65910 105018
rect 65910 104966 65956 105018
rect 65660 104964 65716 104966
rect 65740 104964 65796 104966
rect 65820 104964 65876 104966
rect 65900 104964 65956 104966
rect 65660 103930 65716 103932
rect 65740 103930 65796 103932
rect 65820 103930 65876 103932
rect 65900 103930 65956 103932
rect 65660 103878 65706 103930
rect 65706 103878 65716 103930
rect 65740 103878 65770 103930
rect 65770 103878 65782 103930
rect 65782 103878 65796 103930
rect 65820 103878 65834 103930
rect 65834 103878 65846 103930
rect 65846 103878 65876 103930
rect 65900 103878 65910 103930
rect 65910 103878 65956 103930
rect 65660 103876 65716 103878
rect 65740 103876 65796 103878
rect 65820 103876 65876 103878
rect 65900 103876 65956 103878
rect 65660 102842 65716 102844
rect 65740 102842 65796 102844
rect 65820 102842 65876 102844
rect 65900 102842 65956 102844
rect 65660 102790 65706 102842
rect 65706 102790 65716 102842
rect 65740 102790 65770 102842
rect 65770 102790 65782 102842
rect 65782 102790 65796 102842
rect 65820 102790 65834 102842
rect 65834 102790 65846 102842
rect 65846 102790 65876 102842
rect 65900 102790 65910 102842
rect 65910 102790 65956 102842
rect 65660 102788 65716 102790
rect 65740 102788 65796 102790
rect 65820 102788 65876 102790
rect 65900 102788 65956 102790
rect 65660 101754 65716 101756
rect 65740 101754 65796 101756
rect 65820 101754 65876 101756
rect 65900 101754 65956 101756
rect 65660 101702 65706 101754
rect 65706 101702 65716 101754
rect 65740 101702 65770 101754
rect 65770 101702 65782 101754
rect 65782 101702 65796 101754
rect 65820 101702 65834 101754
rect 65834 101702 65846 101754
rect 65846 101702 65876 101754
rect 65900 101702 65910 101754
rect 65910 101702 65956 101754
rect 65660 101700 65716 101702
rect 65740 101700 65796 101702
rect 65820 101700 65876 101702
rect 65900 101700 65956 101702
rect 65660 100666 65716 100668
rect 65740 100666 65796 100668
rect 65820 100666 65876 100668
rect 65900 100666 65956 100668
rect 65660 100614 65706 100666
rect 65706 100614 65716 100666
rect 65740 100614 65770 100666
rect 65770 100614 65782 100666
rect 65782 100614 65796 100666
rect 65820 100614 65834 100666
rect 65834 100614 65846 100666
rect 65846 100614 65876 100666
rect 65900 100614 65910 100666
rect 65910 100614 65956 100666
rect 65660 100612 65716 100614
rect 65740 100612 65796 100614
rect 65820 100612 65876 100614
rect 65900 100612 65956 100614
rect 65660 99578 65716 99580
rect 65740 99578 65796 99580
rect 65820 99578 65876 99580
rect 65900 99578 65956 99580
rect 65660 99526 65706 99578
rect 65706 99526 65716 99578
rect 65740 99526 65770 99578
rect 65770 99526 65782 99578
rect 65782 99526 65796 99578
rect 65820 99526 65834 99578
rect 65834 99526 65846 99578
rect 65846 99526 65876 99578
rect 65900 99526 65910 99578
rect 65910 99526 65956 99578
rect 65660 99524 65716 99526
rect 65740 99524 65796 99526
rect 65820 99524 65876 99526
rect 65900 99524 65956 99526
rect 65660 98490 65716 98492
rect 65740 98490 65796 98492
rect 65820 98490 65876 98492
rect 65900 98490 65956 98492
rect 65660 98438 65706 98490
rect 65706 98438 65716 98490
rect 65740 98438 65770 98490
rect 65770 98438 65782 98490
rect 65782 98438 65796 98490
rect 65820 98438 65834 98490
rect 65834 98438 65846 98490
rect 65846 98438 65876 98490
rect 65900 98438 65910 98490
rect 65910 98438 65956 98490
rect 65660 98436 65716 98438
rect 65740 98436 65796 98438
rect 65820 98436 65876 98438
rect 65900 98436 65956 98438
rect 65660 97402 65716 97404
rect 65740 97402 65796 97404
rect 65820 97402 65876 97404
rect 65900 97402 65956 97404
rect 65660 97350 65706 97402
rect 65706 97350 65716 97402
rect 65740 97350 65770 97402
rect 65770 97350 65782 97402
rect 65782 97350 65796 97402
rect 65820 97350 65834 97402
rect 65834 97350 65846 97402
rect 65846 97350 65876 97402
rect 65900 97350 65910 97402
rect 65910 97350 65956 97402
rect 65660 97348 65716 97350
rect 65740 97348 65796 97350
rect 65820 97348 65876 97350
rect 65900 97348 65956 97350
rect 65660 96314 65716 96316
rect 65740 96314 65796 96316
rect 65820 96314 65876 96316
rect 65900 96314 65956 96316
rect 65660 96262 65706 96314
rect 65706 96262 65716 96314
rect 65740 96262 65770 96314
rect 65770 96262 65782 96314
rect 65782 96262 65796 96314
rect 65820 96262 65834 96314
rect 65834 96262 65846 96314
rect 65846 96262 65876 96314
rect 65900 96262 65910 96314
rect 65910 96262 65956 96314
rect 65660 96260 65716 96262
rect 65740 96260 65796 96262
rect 65820 96260 65876 96262
rect 65900 96260 65956 96262
rect 65660 95226 65716 95228
rect 65740 95226 65796 95228
rect 65820 95226 65876 95228
rect 65900 95226 65956 95228
rect 65660 95174 65706 95226
rect 65706 95174 65716 95226
rect 65740 95174 65770 95226
rect 65770 95174 65782 95226
rect 65782 95174 65796 95226
rect 65820 95174 65834 95226
rect 65834 95174 65846 95226
rect 65846 95174 65876 95226
rect 65900 95174 65910 95226
rect 65910 95174 65956 95226
rect 65660 95172 65716 95174
rect 65740 95172 65796 95174
rect 65820 95172 65876 95174
rect 65900 95172 65956 95174
rect 65660 94138 65716 94140
rect 65740 94138 65796 94140
rect 65820 94138 65876 94140
rect 65900 94138 65956 94140
rect 65660 94086 65706 94138
rect 65706 94086 65716 94138
rect 65740 94086 65770 94138
rect 65770 94086 65782 94138
rect 65782 94086 65796 94138
rect 65820 94086 65834 94138
rect 65834 94086 65846 94138
rect 65846 94086 65876 94138
rect 65900 94086 65910 94138
rect 65910 94086 65956 94138
rect 65660 94084 65716 94086
rect 65740 94084 65796 94086
rect 65820 94084 65876 94086
rect 65900 94084 65956 94086
rect 65660 93050 65716 93052
rect 65740 93050 65796 93052
rect 65820 93050 65876 93052
rect 65900 93050 65956 93052
rect 65660 92998 65706 93050
rect 65706 92998 65716 93050
rect 65740 92998 65770 93050
rect 65770 92998 65782 93050
rect 65782 92998 65796 93050
rect 65820 92998 65834 93050
rect 65834 92998 65846 93050
rect 65846 92998 65876 93050
rect 65900 92998 65910 93050
rect 65910 92998 65956 93050
rect 65660 92996 65716 92998
rect 65740 92996 65796 92998
rect 65820 92996 65876 92998
rect 65900 92996 65956 92998
rect 65660 91962 65716 91964
rect 65740 91962 65796 91964
rect 65820 91962 65876 91964
rect 65900 91962 65956 91964
rect 65660 91910 65706 91962
rect 65706 91910 65716 91962
rect 65740 91910 65770 91962
rect 65770 91910 65782 91962
rect 65782 91910 65796 91962
rect 65820 91910 65834 91962
rect 65834 91910 65846 91962
rect 65846 91910 65876 91962
rect 65900 91910 65910 91962
rect 65910 91910 65956 91962
rect 65660 91908 65716 91910
rect 65740 91908 65796 91910
rect 65820 91908 65876 91910
rect 65900 91908 65956 91910
rect 65660 90874 65716 90876
rect 65740 90874 65796 90876
rect 65820 90874 65876 90876
rect 65900 90874 65956 90876
rect 65660 90822 65706 90874
rect 65706 90822 65716 90874
rect 65740 90822 65770 90874
rect 65770 90822 65782 90874
rect 65782 90822 65796 90874
rect 65820 90822 65834 90874
rect 65834 90822 65846 90874
rect 65846 90822 65876 90874
rect 65900 90822 65910 90874
rect 65910 90822 65956 90874
rect 65660 90820 65716 90822
rect 65740 90820 65796 90822
rect 65820 90820 65876 90822
rect 65900 90820 65956 90822
rect 65660 89786 65716 89788
rect 65740 89786 65796 89788
rect 65820 89786 65876 89788
rect 65900 89786 65956 89788
rect 65660 89734 65706 89786
rect 65706 89734 65716 89786
rect 65740 89734 65770 89786
rect 65770 89734 65782 89786
rect 65782 89734 65796 89786
rect 65820 89734 65834 89786
rect 65834 89734 65846 89786
rect 65846 89734 65876 89786
rect 65900 89734 65910 89786
rect 65910 89734 65956 89786
rect 65660 89732 65716 89734
rect 65740 89732 65796 89734
rect 65820 89732 65876 89734
rect 65900 89732 65956 89734
rect 65660 88698 65716 88700
rect 65740 88698 65796 88700
rect 65820 88698 65876 88700
rect 65900 88698 65956 88700
rect 65660 88646 65706 88698
rect 65706 88646 65716 88698
rect 65740 88646 65770 88698
rect 65770 88646 65782 88698
rect 65782 88646 65796 88698
rect 65820 88646 65834 88698
rect 65834 88646 65846 88698
rect 65846 88646 65876 88698
rect 65900 88646 65910 88698
rect 65910 88646 65956 88698
rect 65660 88644 65716 88646
rect 65740 88644 65796 88646
rect 65820 88644 65876 88646
rect 65900 88644 65956 88646
rect 65660 87610 65716 87612
rect 65740 87610 65796 87612
rect 65820 87610 65876 87612
rect 65900 87610 65956 87612
rect 65660 87558 65706 87610
rect 65706 87558 65716 87610
rect 65740 87558 65770 87610
rect 65770 87558 65782 87610
rect 65782 87558 65796 87610
rect 65820 87558 65834 87610
rect 65834 87558 65846 87610
rect 65846 87558 65876 87610
rect 65900 87558 65910 87610
rect 65910 87558 65956 87610
rect 65660 87556 65716 87558
rect 65740 87556 65796 87558
rect 65820 87556 65876 87558
rect 65900 87556 65956 87558
rect 65660 86522 65716 86524
rect 65740 86522 65796 86524
rect 65820 86522 65876 86524
rect 65900 86522 65956 86524
rect 65660 86470 65706 86522
rect 65706 86470 65716 86522
rect 65740 86470 65770 86522
rect 65770 86470 65782 86522
rect 65782 86470 65796 86522
rect 65820 86470 65834 86522
rect 65834 86470 65846 86522
rect 65846 86470 65876 86522
rect 65900 86470 65910 86522
rect 65910 86470 65956 86522
rect 65660 86468 65716 86470
rect 65740 86468 65796 86470
rect 65820 86468 65876 86470
rect 65900 86468 65956 86470
rect 65660 85434 65716 85436
rect 65740 85434 65796 85436
rect 65820 85434 65876 85436
rect 65900 85434 65956 85436
rect 65660 85382 65706 85434
rect 65706 85382 65716 85434
rect 65740 85382 65770 85434
rect 65770 85382 65782 85434
rect 65782 85382 65796 85434
rect 65820 85382 65834 85434
rect 65834 85382 65846 85434
rect 65846 85382 65876 85434
rect 65900 85382 65910 85434
rect 65910 85382 65956 85434
rect 65660 85380 65716 85382
rect 65740 85380 65796 85382
rect 65820 85380 65876 85382
rect 65900 85380 65956 85382
rect 65660 84346 65716 84348
rect 65740 84346 65796 84348
rect 65820 84346 65876 84348
rect 65900 84346 65956 84348
rect 65660 84294 65706 84346
rect 65706 84294 65716 84346
rect 65740 84294 65770 84346
rect 65770 84294 65782 84346
rect 65782 84294 65796 84346
rect 65820 84294 65834 84346
rect 65834 84294 65846 84346
rect 65846 84294 65876 84346
rect 65900 84294 65910 84346
rect 65910 84294 65956 84346
rect 65660 84292 65716 84294
rect 65740 84292 65796 84294
rect 65820 84292 65876 84294
rect 65900 84292 65956 84294
rect 65660 83258 65716 83260
rect 65740 83258 65796 83260
rect 65820 83258 65876 83260
rect 65900 83258 65956 83260
rect 65660 83206 65706 83258
rect 65706 83206 65716 83258
rect 65740 83206 65770 83258
rect 65770 83206 65782 83258
rect 65782 83206 65796 83258
rect 65820 83206 65834 83258
rect 65834 83206 65846 83258
rect 65846 83206 65876 83258
rect 65900 83206 65910 83258
rect 65910 83206 65956 83258
rect 65660 83204 65716 83206
rect 65740 83204 65796 83206
rect 65820 83204 65876 83206
rect 65900 83204 65956 83206
rect 65660 82170 65716 82172
rect 65740 82170 65796 82172
rect 65820 82170 65876 82172
rect 65900 82170 65956 82172
rect 65660 82118 65706 82170
rect 65706 82118 65716 82170
rect 65740 82118 65770 82170
rect 65770 82118 65782 82170
rect 65782 82118 65796 82170
rect 65820 82118 65834 82170
rect 65834 82118 65846 82170
rect 65846 82118 65876 82170
rect 65900 82118 65910 82170
rect 65910 82118 65956 82170
rect 65660 82116 65716 82118
rect 65740 82116 65796 82118
rect 65820 82116 65876 82118
rect 65900 82116 65956 82118
rect 65660 81082 65716 81084
rect 65740 81082 65796 81084
rect 65820 81082 65876 81084
rect 65900 81082 65956 81084
rect 65660 81030 65706 81082
rect 65706 81030 65716 81082
rect 65740 81030 65770 81082
rect 65770 81030 65782 81082
rect 65782 81030 65796 81082
rect 65820 81030 65834 81082
rect 65834 81030 65846 81082
rect 65846 81030 65876 81082
rect 65900 81030 65910 81082
rect 65910 81030 65956 81082
rect 65660 81028 65716 81030
rect 65740 81028 65796 81030
rect 65820 81028 65876 81030
rect 65900 81028 65956 81030
rect 65660 79994 65716 79996
rect 65740 79994 65796 79996
rect 65820 79994 65876 79996
rect 65900 79994 65956 79996
rect 65660 79942 65706 79994
rect 65706 79942 65716 79994
rect 65740 79942 65770 79994
rect 65770 79942 65782 79994
rect 65782 79942 65796 79994
rect 65820 79942 65834 79994
rect 65834 79942 65846 79994
rect 65846 79942 65876 79994
rect 65900 79942 65910 79994
rect 65910 79942 65956 79994
rect 65660 79940 65716 79942
rect 65740 79940 65796 79942
rect 65820 79940 65876 79942
rect 65900 79940 65956 79942
rect 65660 78906 65716 78908
rect 65740 78906 65796 78908
rect 65820 78906 65876 78908
rect 65900 78906 65956 78908
rect 65660 78854 65706 78906
rect 65706 78854 65716 78906
rect 65740 78854 65770 78906
rect 65770 78854 65782 78906
rect 65782 78854 65796 78906
rect 65820 78854 65834 78906
rect 65834 78854 65846 78906
rect 65846 78854 65876 78906
rect 65900 78854 65910 78906
rect 65910 78854 65956 78906
rect 65660 78852 65716 78854
rect 65740 78852 65796 78854
rect 65820 78852 65876 78854
rect 65900 78852 65956 78854
rect 65660 77818 65716 77820
rect 65740 77818 65796 77820
rect 65820 77818 65876 77820
rect 65900 77818 65956 77820
rect 65660 77766 65706 77818
rect 65706 77766 65716 77818
rect 65740 77766 65770 77818
rect 65770 77766 65782 77818
rect 65782 77766 65796 77818
rect 65820 77766 65834 77818
rect 65834 77766 65846 77818
rect 65846 77766 65876 77818
rect 65900 77766 65910 77818
rect 65910 77766 65956 77818
rect 65660 77764 65716 77766
rect 65740 77764 65796 77766
rect 65820 77764 65876 77766
rect 65900 77764 65956 77766
rect 65660 76730 65716 76732
rect 65740 76730 65796 76732
rect 65820 76730 65876 76732
rect 65900 76730 65956 76732
rect 65660 76678 65706 76730
rect 65706 76678 65716 76730
rect 65740 76678 65770 76730
rect 65770 76678 65782 76730
rect 65782 76678 65796 76730
rect 65820 76678 65834 76730
rect 65834 76678 65846 76730
rect 65846 76678 65876 76730
rect 65900 76678 65910 76730
rect 65910 76678 65956 76730
rect 65660 76676 65716 76678
rect 65740 76676 65796 76678
rect 65820 76676 65876 76678
rect 65900 76676 65956 76678
rect 65660 75642 65716 75644
rect 65740 75642 65796 75644
rect 65820 75642 65876 75644
rect 65900 75642 65956 75644
rect 65660 75590 65706 75642
rect 65706 75590 65716 75642
rect 65740 75590 65770 75642
rect 65770 75590 65782 75642
rect 65782 75590 65796 75642
rect 65820 75590 65834 75642
rect 65834 75590 65846 75642
rect 65846 75590 65876 75642
rect 65900 75590 65910 75642
rect 65910 75590 65956 75642
rect 65660 75588 65716 75590
rect 65740 75588 65796 75590
rect 65820 75588 65876 75590
rect 65900 75588 65956 75590
rect 65660 74554 65716 74556
rect 65740 74554 65796 74556
rect 65820 74554 65876 74556
rect 65900 74554 65956 74556
rect 65660 74502 65706 74554
rect 65706 74502 65716 74554
rect 65740 74502 65770 74554
rect 65770 74502 65782 74554
rect 65782 74502 65796 74554
rect 65820 74502 65834 74554
rect 65834 74502 65846 74554
rect 65846 74502 65876 74554
rect 65900 74502 65910 74554
rect 65910 74502 65956 74554
rect 65660 74500 65716 74502
rect 65740 74500 65796 74502
rect 65820 74500 65876 74502
rect 65900 74500 65956 74502
rect 65660 73466 65716 73468
rect 65740 73466 65796 73468
rect 65820 73466 65876 73468
rect 65900 73466 65956 73468
rect 65660 73414 65706 73466
rect 65706 73414 65716 73466
rect 65740 73414 65770 73466
rect 65770 73414 65782 73466
rect 65782 73414 65796 73466
rect 65820 73414 65834 73466
rect 65834 73414 65846 73466
rect 65846 73414 65876 73466
rect 65900 73414 65910 73466
rect 65910 73414 65956 73466
rect 65660 73412 65716 73414
rect 65740 73412 65796 73414
rect 65820 73412 65876 73414
rect 65900 73412 65956 73414
rect 65660 72378 65716 72380
rect 65740 72378 65796 72380
rect 65820 72378 65876 72380
rect 65900 72378 65956 72380
rect 65660 72326 65706 72378
rect 65706 72326 65716 72378
rect 65740 72326 65770 72378
rect 65770 72326 65782 72378
rect 65782 72326 65796 72378
rect 65820 72326 65834 72378
rect 65834 72326 65846 72378
rect 65846 72326 65876 72378
rect 65900 72326 65910 72378
rect 65910 72326 65956 72378
rect 65660 72324 65716 72326
rect 65740 72324 65796 72326
rect 65820 72324 65876 72326
rect 65900 72324 65956 72326
rect 65660 71290 65716 71292
rect 65740 71290 65796 71292
rect 65820 71290 65876 71292
rect 65900 71290 65956 71292
rect 65660 71238 65706 71290
rect 65706 71238 65716 71290
rect 65740 71238 65770 71290
rect 65770 71238 65782 71290
rect 65782 71238 65796 71290
rect 65820 71238 65834 71290
rect 65834 71238 65846 71290
rect 65846 71238 65876 71290
rect 65900 71238 65910 71290
rect 65910 71238 65956 71290
rect 65660 71236 65716 71238
rect 65740 71236 65796 71238
rect 65820 71236 65876 71238
rect 65900 71236 65956 71238
rect 65660 70202 65716 70204
rect 65740 70202 65796 70204
rect 65820 70202 65876 70204
rect 65900 70202 65956 70204
rect 65660 70150 65706 70202
rect 65706 70150 65716 70202
rect 65740 70150 65770 70202
rect 65770 70150 65782 70202
rect 65782 70150 65796 70202
rect 65820 70150 65834 70202
rect 65834 70150 65846 70202
rect 65846 70150 65876 70202
rect 65900 70150 65910 70202
rect 65910 70150 65956 70202
rect 65660 70148 65716 70150
rect 65740 70148 65796 70150
rect 65820 70148 65876 70150
rect 65900 70148 65956 70150
rect 65660 69114 65716 69116
rect 65740 69114 65796 69116
rect 65820 69114 65876 69116
rect 65900 69114 65956 69116
rect 65660 69062 65706 69114
rect 65706 69062 65716 69114
rect 65740 69062 65770 69114
rect 65770 69062 65782 69114
rect 65782 69062 65796 69114
rect 65820 69062 65834 69114
rect 65834 69062 65846 69114
rect 65846 69062 65876 69114
rect 65900 69062 65910 69114
rect 65910 69062 65956 69114
rect 65660 69060 65716 69062
rect 65740 69060 65796 69062
rect 65820 69060 65876 69062
rect 65900 69060 65956 69062
rect 65660 68026 65716 68028
rect 65740 68026 65796 68028
rect 65820 68026 65876 68028
rect 65900 68026 65956 68028
rect 65660 67974 65706 68026
rect 65706 67974 65716 68026
rect 65740 67974 65770 68026
rect 65770 67974 65782 68026
rect 65782 67974 65796 68026
rect 65820 67974 65834 68026
rect 65834 67974 65846 68026
rect 65846 67974 65876 68026
rect 65900 67974 65910 68026
rect 65910 67974 65956 68026
rect 65660 67972 65716 67974
rect 65740 67972 65796 67974
rect 65820 67972 65876 67974
rect 65900 67972 65956 67974
rect 65660 66938 65716 66940
rect 65740 66938 65796 66940
rect 65820 66938 65876 66940
rect 65900 66938 65956 66940
rect 65660 66886 65706 66938
rect 65706 66886 65716 66938
rect 65740 66886 65770 66938
rect 65770 66886 65782 66938
rect 65782 66886 65796 66938
rect 65820 66886 65834 66938
rect 65834 66886 65846 66938
rect 65846 66886 65876 66938
rect 65900 66886 65910 66938
rect 65910 66886 65956 66938
rect 65660 66884 65716 66886
rect 65740 66884 65796 66886
rect 65820 66884 65876 66886
rect 65900 66884 65956 66886
rect 65660 65850 65716 65852
rect 65740 65850 65796 65852
rect 65820 65850 65876 65852
rect 65900 65850 65956 65852
rect 65660 65798 65706 65850
rect 65706 65798 65716 65850
rect 65740 65798 65770 65850
rect 65770 65798 65782 65850
rect 65782 65798 65796 65850
rect 65820 65798 65834 65850
rect 65834 65798 65846 65850
rect 65846 65798 65876 65850
rect 65900 65798 65910 65850
rect 65910 65798 65956 65850
rect 65660 65796 65716 65798
rect 65740 65796 65796 65798
rect 65820 65796 65876 65798
rect 65900 65796 65956 65798
rect 65660 64762 65716 64764
rect 65740 64762 65796 64764
rect 65820 64762 65876 64764
rect 65900 64762 65956 64764
rect 65660 64710 65706 64762
rect 65706 64710 65716 64762
rect 65740 64710 65770 64762
rect 65770 64710 65782 64762
rect 65782 64710 65796 64762
rect 65820 64710 65834 64762
rect 65834 64710 65846 64762
rect 65846 64710 65876 64762
rect 65900 64710 65910 64762
rect 65910 64710 65956 64762
rect 65660 64708 65716 64710
rect 65740 64708 65796 64710
rect 65820 64708 65876 64710
rect 65900 64708 65956 64710
rect 65660 63674 65716 63676
rect 65740 63674 65796 63676
rect 65820 63674 65876 63676
rect 65900 63674 65956 63676
rect 65660 63622 65706 63674
rect 65706 63622 65716 63674
rect 65740 63622 65770 63674
rect 65770 63622 65782 63674
rect 65782 63622 65796 63674
rect 65820 63622 65834 63674
rect 65834 63622 65846 63674
rect 65846 63622 65876 63674
rect 65900 63622 65910 63674
rect 65910 63622 65956 63674
rect 65660 63620 65716 63622
rect 65740 63620 65796 63622
rect 65820 63620 65876 63622
rect 65900 63620 65956 63622
rect 65660 62586 65716 62588
rect 65740 62586 65796 62588
rect 65820 62586 65876 62588
rect 65900 62586 65956 62588
rect 65660 62534 65706 62586
rect 65706 62534 65716 62586
rect 65740 62534 65770 62586
rect 65770 62534 65782 62586
rect 65782 62534 65796 62586
rect 65820 62534 65834 62586
rect 65834 62534 65846 62586
rect 65846 62534 65876 62586
rect 65900 62534 65910 62586
rect 65910 62534 65956 62586
rect 65660 62532 65716 62534
rect 65740 62532 65796 62534
rect 65820 62532 65876 62534
rect 65900 62532 65956 62534
rect 65660 61498 65716 61500
rect 65740 61498 65796 61500
rect 65820 61498 65876 61500
rect 65900 61498 65956 61500
rect 65660 61446 65706 61498
rect 65706 61446 65716 61498
rect 65740 61446 65770 61498
rect 65770 61446 65782 61498
rect 65782 61446 65796 61498
rect 65820 61446 65834 61498
rect 65834 61446 65846 61498
rect 65846 61446 65876 61498
rect 65900 61446 65910 61498
rect 65910 61446 65956 61498
rect 65660 61444 65716 61446
rect 65740 61444 65796 61446
rect 65820 61444 65876 61446
rect 65900 61444 65956 61446
rect 65660 60410 65716 60412
rect 65740 60410 65796 60412
rect 65820 60410 65876 60412
rect 65900 60410 65956 60412
rect 65660 60358 65706 60410
rect 65706 60358 65716 60410
rect 65740 60358 65770 60410
rect 65770 60358 65782 60410
rect 65782 60358 65796 60410
rect 65820 60358 65834 60410
rect 65834 60358 65846 60410
rect 65846 60358 65876 60410
rect 65900 60358 65910 60410
rect 65910 60358 65956 60410
rect 65660 60356 65716 60358
rect 65740 60356 65796 60358
rect 65820 60356 65876 60358
rect 65900 60356 65956 60358
rect 78034 114316 78036 114336
rect 78036 114316 78088 114336
rect 78088 114316 78090 114336
rect 78034 114280 78090 114316
rect 77574 78920 77630 78976
rect 65660 59322 65716 59324
rect 65740 59322 65796 59324
rect 65820 59322 65876 59324
rect 65900 59322 65956 59324
rect 65660 59270 65706 59322
rect 65706 59270 65716 59322
rect 65740 59270 65770 59322
rect 65770 59270 65782 59322
rect 65782 59270 65796 59322
rect 65820 59270 65834 59322
rect 65834 59270 65846 59322
rect 65846 59270 65876 59322
rect 65900 59270 65910 59322
rect 65910 59270 65956 59322
rect 65660 59268 65716 59270
rect 65740 59268 65796 59270
rect 65820 59268 65876 59270
rect 65900 59268 65956 59270
rect 65660 58234 65716 58236
rect 65740 58234 65796 58236
rect 65820 58234 65876 58236
rect 65900 58234 65956 58236
rect 65660 58182 65706 58234
rect 65706 58182 65716 58234
rect 65740 58182 65770 58234
rect 65770 58182 65782 58234
rect 65782 58182 65796 58234
rect 65820 58182 65834 58234
rect 65834 58182 65846 58234
rect 65846 58182 65876 58234
rect 65900 58182 65910 58234
rect 65910 58182 65956 58234
rect 65660 58180 65716 58182
rect 65740 58180 65796 58182
rect 65820 58180 65876 58182
rect 65900 58180 65956 58182
rect 65660 57146 65716 57148
rect 65740 57146 65796 57148
rect 65820 57146 65876 57148
rect 65900 57146 65956 57148
rect 65660 57094 65706 57146
rect 65706 57094 65716 57146
rect 65740 57094 65770 57146
rect 65770 57094 65782 57146
rect 65782 57094 65796 57146
rect 65820 57094 65834 57146
rect 65834 57094 65846 57146
rect 65846 57094 65876 57146
rect 65900 57094 65910 57146
rect 65910 57094 65956 57146
rect 65660 57092 65716 57094
rect 65740 57092 65796 57094
rect 65820 57092 65876 57094
rect 65900 57092 65956 57094
rect 65660 56058 65716 56060
rect 65740 56058 65796 56060
rect 65820 56058 65876 56060
rect 65900 56058 65956 56060
rect 65660 56006 65706 56058
rect 65706 56006 65716 56058
rect 65740 56006 65770 56058
rect 65770 56006 65782 56058
rect 65782 56006 65796 56058
rect 65820 56006 65834 56058
rect 65834 56006 65846 56058
rect 65846 56006 65876 56058
rect 65900 56006 65910 56058
rect 65910 56006 65956 56058
rect 65660 56004 65716 56006
rect 65740 56004 65796 56006
rect 65820 56004 65876 56006
rect 65900 56004 65956 56006
rect 65660 54970 65716 54972
rect 65740 54970 65796 54972
rect 65820 54970 65876 54972
rect 65900 54970 65956 54972
rect 65660 54918 65706 54970
rect 65706 54918 65716 54970
rect 65740 54918 65770 54970
rect 65770 54918 65782 54970
rect 65782 54918 65796 54970
rect 65820 54918 65834 54970
rect 65834 54918 65846 54970
rect 65846 54918 65876 54970
rect 65900 54918 65910 54970
rect 65910 54918 65956 54970
rect 65660 54916 65716 54918
rect 65740 54916 65796 54918
rect 65820 54916 65876 54918
rect 65900 54916 65956 54918
rect 65660 53882 65716 53884
rect 65740 53882 65796 53884
rect 65820 53882 65876 53884
rect 65900 53882 65956 53884
rect 65660 53830 65706 53882
rect 65706 53830 65716 53882
rect 65740 53830 65770 53882
rect 65770 53830 65782 53882
rect 65782 53830 65796 53882
rect 65820 53830 65834 53882
rect 65834 53830 65846 53882
rect 65846 53830 65876 53882
rect 65900 53830 65910 53882
rect 65910 53830 65956 53882
rect 65660 53828 65716 53830
rect 65740 53828 65796 53830
rect 65820 53828 65876 53830
rect 65900 53828 65956 53830
rect 65660 52794 65716 52796
rect 65740 52794 65796 52796
rect 65820 52794 65876 52796
rect 65900 52794 65956 52796
rect 65660 52742 65706 52794
rect 65706 52742 65716 52794
rect 65740 52742 65770 52794
rect 65770 52742 65782 52794
rect 65782 52742 65796 52794
rect 65820 52742 65834 52794
rect 65834 52742 65846 52794
rect 65846 52742 65876 52794
rect 65900 52742 65910 52794
rect 65910 52742 65956 52794
rect 65660 52740 65716 52742
rect 65740 52740 65796 52742
rect 65820 52740 65876 52742
rect 65900 52740 65956 52742
rect 65660 51706 65716 51708
rect 65740 51706 65796 51708
rect 65820 51706 65876 51708
rect 65900 51706 65956 51708
rect 65660 51654 65706 51706
rect 65706 51654 65716 51706
rect 65740 51654 65770 51706
rect 65770 51654 65782 51706
rect 65782 51654 65796 51706
rect 65820 51654 65834 51706
rect 65834 51654 65846 51706
rect 65846 51654 65876 51706
rect 65900 51654 65910 51706
rect 65910 51654 65956 51706
rect 65660 51652 65716 51654
rect 65740 51652 65796 51654
rect 65820 51652 65876 51654
rect 65900 51652 65956 51654
rect 65660 50618 65716 50620
rect 65740 50618 65796 50620
rect 65820 50618 65876 50620
rect 65900 50618 65956 50620
rect 65660 50566 65706 50618
rect 65706 50566 65716 50618
rect 65740 50566 65770 50618
rect 65770 50566 65782 50618
rect 65782 50566 65796 50618
rect 65820 50566 65834 50618
rect 65834 50566 65846 50618
rect 65846 50566 65876 50618
rect 65900 50566 65910 50618
rect 65910 50566 65956 50618
rect 65660 50564 65716 50566
rect 65740 50564 65796 50566
rect 65820 50564 65876 50566
rect 65900 50564 65956 50566
rect 65660 49530 65716 49532
rect 65740 49530 65796 49532
rect 65820 49530 65876 49532
rect 65900 49530 65956 49532
rect 65660 49478 65706 49530
rect 65706 49478 65716 49530
rect 65740 49478 65770 49530
rect 65770 49478 65782 49530
rect 65782 49478 65796 49530
rect 65820 49478 65834 49530
rect 65834 49478 65846 49530
rect 65846 49478 65876 49530
rect 65900 49478 65910 49530
rect 65910 49478 65956 49530
rect 65660 49476 65716 49478
rect 65740 49476 65796 49478
rect 65820 49476 65876 49478
rect 65900 49476 65956 49478
rect 65660 48442 65716 48444
rect 65740 48442 65796 48444
rect 65820 48442 65876 48444
rect 65900 48442 65956 48444
rect 65660 48390 65706 48442
rect 65706 48390 65716 48442
rect 65740 48390 65770 48442
rect 65770 48390 65782 48442
rect 65782 48390 65796 48442
rect 65820 48390 65834 48442
rect 65834 48390 65846 48442
rect 65846 48390 65876 48442
rect 65900 48390 65910 48442
rect 65910 48390 65956 48442
rect 65660 48388 65716 48390
rect 65740 48388 65796 48390
rect 65820 48388 65876 48390
rect 65900 48388 65956 48390
rect 75826 47640 75882 47696
rect 65660 47354 65716 47356
rect 65740 47354 65796 47356
rect 65820 47354 65876 47356
rect 65900 47354 65956 47356
rect 65660 47302 65706 47354
rect 65706 47302 65716 47354
rect 65740 47302 65770 47354
rect 65770 47302 65782 47354
rect 65782 47302 65796 47354
rect 65820 47302 65834 47354
rect 65834 47302 65846 47354
rect 65846 47302 65876 47354
rect 65900 47302 65910 47354
rect 65910 47302 65956 47354
rect 65660 47300 65716 47302
rect 65740 47300 65796 47302
rect 65820 47300 65876 47302
rect 65900 47300 65956 47302
rect 65660 46266 65716 46268
rect 65740 46266 65796 46268
rect 65820 46266 65876 46268
rect 65900 46266 65956 46268
rect 65660 46214 65706 46266
rect 65706 46214 65716 46266
rect 65740 46214 65770 46266
rect 65770 46214 65782 46266
rect 65782 46214 65796 46266
rect 65820 46214 65834 46266
rect 65834 46214 65846 46266
rect 65846 46214 65876 46266
rect 65900 46214 65910 46266
rect 65910 46214 65956 46266
rect 65660 46212 65716 46214
rect 65740 46212 65796 46214
rect 65820 46212 65876 46214
rect 65900 46212 65956 46214
rect 65660 45178 65716 45180
rect 65740 45178 65796 45180
rect 65820 45178 65876 45180
rect 65900 45178 65956 45180
rect 65660 45126 65706 45178
rect 65706 45126 65716 45178
rect 65740 45126 65770 45178
rect 65770 45126 65782 45178
rect 65782 45126 65796 45178
rect 65820 45126 65834 45178
rect 65834 45126 65846 45178
rect 65846 45126 65876 45178
rect 65900 45126 65910 45178
rect 65910 45126 65956 45178
rect 65660 45124 65716 45126
rect 65740 45124 65796 45126
rect 65820 45124 65876 45126
rect 65900 45124 65956 45126
rect 65660 44090 65716 44092
rect 65740 44090 65796 44092
rect 65820 44090 65876 44092
rect 65900 44090 65956 44092
rect 65660 44038 65706 44090
rect 65706 44038 65716 44090
rect 65740 44038 65770 44090
rect 65770 44038 65782 44090
rect 65782 44038 65796 44090
rect 65820 44038 65834 44090
rect 65834 44038 65846 44090
rect 65846 44038 65876 44090
rect 65900 44038 65910 44090
rect 65910 44038 65956 44090
rect 65660 44036 65716 44038
rect 65740 44036 65796 44038
rect 65820 44036 65876 44038
rect 65900 44036 65956 44038
rect 65660 43002 65716 43004
rect 65740 43002 65796 43004
rect 65820 43002 65876 43004
rect 65900 43002 65956 43004
rect 65660 42950 65706 43002
rect 65706 42950 65716 43002
rect 65740 42950 65770 43002
rect 65770 42950 65782 43002
rect 65782 42950 65796 43002
rect 65820 42950 65834 43002
rect 65834 42950 65846 43002
rect 65846 42950 65876 43002
rect 65900 42950 65910 43002
rect 65910 42950 65956 43002
rect 65660 42948 65716 42950
rect 65740 42948 65796 42950
rect 65820 42948 65876 42950
rect 65900 42948 65956 42950
rect 65660 41914 65716 41916
rect 65740 41914 65796 41916
rect 65820 41914 65876 41916
rect 65900 41914 65956 41916
rect 65660 41862 65706 41914
rect 65706 41862 65716 41914
rect 65740 41862 65770 41914
rect 65770 41862 65782 41914
rect 65782 41862 65796 41914
rect 65820 41862 65834 41914
rect 65834 41862 65846 41914
rect 65846 41862 65876 41914
rect 65900 41862 65910 41914
rect 65910 41862 65956 41914
rect 65660 41860 65716 41862
rect 65740 41860 65796 41862
rect 65820 41860 65876 41862
rect 65900 41860 65956 41862
rect 65660 40826 65716 40828
rect 65740 40826 65796 40828
rect 65820 40826 65876 40828
rect 65900 40826 65956 40828
rect 65660 40774 65706 40826
rect 65706 40774 65716 40826
rect 65740 40774 65770 40826
rect 65770 40774 65782 40826
rect 65782 40774 65796 40826
rect 65820 40774 65834 40826
rect 65834 40774 65846 40826
rect 65846 40774 65876 40826
rect 65900 40774 65910 40826
rect 65910 40774 65956 40826
rect 65660 40772 65716 40774
rect 65740 40772 65796 40774
rect 65820 40772 65876 40774
rect 65900 40772 65956 40774
rect 65660 39738 65716 39740
rect 65740 39738 65796 39740
rect 65820 39738 65876 39740
rect 65900 39738 65956 39740
rect 65660 39686 65706 39738
rect 65706 39686 65716 39738
rect 65740 39686 65770 39738
rect 65770 39686 65782 39738
rect 65782 39686 65796 39738
rect 65820 39686 65834 39738
rect 65834 39686 65846 39738
rect 65846 39686 65876 39738
rect 65900 39686 65910 39738
rect 65910 39686 65956 39738
rect 65660 39684 65716 39686
rect 65740 39684 65796 39686
rect 65820 39684 65876 39686
rect 65900 39684 65956 39686
rect 65660 38650 65716 38652
rect 65740 38650 65796 38652
rect 65820 38650 65876 38652
rect 65900 38650 65956 38652
rect 65660 38598 65706 38650
rect 65706 38598 65716 38650
rect 65740 38598 65770 38650
rect 65770 38598 65782 38650
rect 65782 38598 65796 38650
rect 65820 38598 65834 38650
rect 65834 38598 65846 38650
rect 65846 38598 65876 38650
rect 65900 38598 65910 38650
rect 65910 38598 65956 38650
rect 65660 38596 65716 38598
rect 65740 38596 65796 38598
rect 65820 38596 65876 38598
rect 65900 38596 65956 38598
rect 65660 37562 65716 37564
rect 65740 37562 65796 37564
rect 65820 37562 65876 37564
rect 65900 37562 65956 37564
rect 65660 37510 65706 37562
rect 65706 37510 65716 37562
rect 65740 37510 65770 37562
rect 65770 37510 65782 37562
rect 65782 37510 65796 37562
rect 65820 37510 65834 37562
rect 65834 37510 65846 37562
rect 65846 37510 65876 37562
rect 65900 37510 65910 37562
rect 65910 37510 65956 37562
rect 65660 37508 65716 37510
rect 65740 37508 65796 37510
rect 65820 37508 65876 37510
rect 65900 37508 65956 37510
rect 65660 36474 65716 36476
rect 65740 36474 65796 36476
rect 65820 36474 65876 36476
rect 65900 36474 65956 36476
rect 65660 36422 65706 36474
rect 65706 36422 65716 36474
rect 65740 36422 65770 36474
rect 65770 36422 65782 36474
rect 65782 36422 65796 36474
rect 65820 36422 65834 36474
rect 65834 36422 65846 36474
rect 65846 36422 65876 36474
rect 65900 36422 65910 36474
rect 65910 36422 65956 36474
rect 65660 36420 65716 36422
rect 65740 36420 65796 36422
rect 65820 36420 65876 36422
rect 65900 36420 65956 36422
rect 65660 35386 65716 35388
rect 65740 35386 65796 35388
rect 65820 35386 65876 35388
rect 65900 35386 65956 35388
rect 65660 35334 65706 35386
rect 65706 35334 65716 35386
rect 65740 35334 65770 35386
rect 65770 35334 65782 35386
rect 65782 35334 65796 35386
rect 65820 35334 65834 35386
rect 65834 35334 65846 35386
rect 65846 35334 65876 35386
rect 65900 35334 65910 35386
rect 65910 35334 65956 35386
rect 65660 35332 65716 35334
rect 65740 35332 65796 35334
rect 65820 35332 65876 35334
rect 65900 35332 65956 35334
rect 65660 34298 65716 34300
rect 65740 34298 65796 34300
rect 65820 34298 65876 34300
rect 65900 34298 65956 34300
rect 65660 34246 65706 34298
rect 65706 34246 65716 34298
rect 65740 34246 65770 34298
rect 65770 34246 65782 34298
rect 65782 34246 65796 34298
rect 65820 34246 65834 34298
rect 65834 34246 65846 34298
rect 65846 34246 65876 34298
rect 65900 34246 65910 34298
rect 65910 34246 65956 34298
rect 65660 34244 65716 34246
rect 65740 34244 65796 34246
rect 65820 34244 65876 34246
rect 65900 34244 65956 34246
rect 65660 33210 65716 33212
rect 65740 33210 65796 33212
rect 65820 33210 65876 33212
rect 65900 33210 65956 33212
rect 65660 33158 65706 33210
rect 65706 33158 65716 33210
rect 65740 33158 65770 33210
rect 65770 33158 65782 33210
rect 65782 33158 65796 33210
rect 65820 33158 65834 33210
rect 65834 33158 65846 33210
rect 65846 33158 65876 33210
rect 65900 33158 65910 33210
rect 65910 33158 65956 33210
rect 65660 33156 65716 33158
rect 65740 33156 65796 33158
rect 65820 33156 65876 33158
rect 65900 33156 65956 33158
rect 65660 32122 65716 32124
rect 65740 32122 65796 32124
rect 65820 32122 65876 32124
rect 65900 32122 65956 32124
rect 65660 32070 65706 32122
rect 65706 32070 65716 32122
rect 65740 32070 65770 32122
rect 65770 32070 65782 32122
rect 65782 32070 65796 32122
rect 65820 32070 65834 32122
rect 65834 32070 65846 32122
rect 65846 32070 65876 32122
rect 65900 32070 65910 32122
rect 65910 32070 65956 32122
rect 65660 32068 65716 32070
rect 65740 32068 65796 32070
rect 65820 32068 65876 32070
rect 65900 32068 65956 32070
rect 65660 31034 65716 31036
rect 65740 31034 65796 31036
rect 65820 31034 65876 31036
rect 65900 31034 65956 31036
rect 65660 30982 65706 31034
rect 65706 30982 65716 31034
rect 65740 30982 65770 31034
rect 65770 30982 65782 31034
rect 65782 30982 65796 31034
rect 65820 30982 65834 31034
rect 65834 30982 65846 31034
rect 65846 30982 65876 31034
rect 65900 30982 65910 31034
rect 65910 30982 65956 31034
rect 65660 30980 65716 30982
rect 65740 30980 65796 30982
rect 65820 30980 65876 30982
rect 65900 30980 65956 30982
rect 65660 29946 65716 29948
rect 65740 29946 65796 29948
rect 65820 29946 65876 29948
rect 65900 29946 65956 29948
rect 65660 29894 65706 29946
rect 65706 29894 65716 29946
rect 65740 29894 65770 29946
rect 65770 29894 65782 29946
rect 65782 29894 65796 29946
rect 65820 29894 65834 29946
rect 65834 29894 65846 29946
rect 65846 29894 65876 29946
rect 65900 29894 65910 29946
rect 65910 29894 65956 29946
rect 65660 29892 65716 29894
rect 65740 29892 65796 29894
rect 65820 29892 65876 29894
rect 65900 29892 65956 29894
rect 65660 28858 65716 28860
rect 65740 28858 65796 28860
rect 65820 28858 65876 28860
rect 65900 28858 65956 28860
rect 65660 28806 65706 28858
rect 65706 28806 65716 28858
rect 65740 28806 65770 28858
rect 65770 28806 65782 28858
rect 65782 28806 65796 28858
rect 65820 28806 65834 28858
rect 65834 28806 65846 28858
rect 65846 28806 65876 28858
rect 65900 28806 65910 28858
rect 65910 28806 65956 28858
rect 65660 28804 65716 28806
rect 65740 28804 65796 28806
rect 65820 28804 65876 28806
rect 65900 28804 65956 28806
rect 65660 27770 65716 27772
rect 65740 27770 65796 27772
rect 65820 27770 65876 27772
rect 65900 27770 65956 27772
rect 65660 27718 65706 27770
rect 65706 27718 65716 27770
rect 65740 27718 65770 27770
rect 65770 27718 65782 27770
rect 65782 27718 65796 27770
rect 65820 27718 65834 27770
rect 65834 27718 65846 27770
rect 65846 27718 65876 27770
rect 65900 27718 65910 27770
rect 65910 27718 65956 27770
rect 65660 27716 65716 27718
rect 65740 27716 65796 27718
rect 65820 27716 65876 27718
rect 65900 27716 65956 27718
rect 65660 26682 65716 26684
rect 65740 26682 65796 26684
rect 65820 26682 65876 26684
rect 65900 26682 65956 26684
rect 65660 26630 65706 26682
rect 65706 26630 65716 26682
rect 65740 26630 65770 26682
rect 65770 26630 65782 26682
rect 65782 26630 65796 26682
rect 65820 26630 65834 26682
rect 65834 26630 65846 26682
rect 65846 26630 65876 26682
rect 65900 26630 65910 26682
rect 65910 26630 65956 26682
rect 65660 26628 65716 26630
rect 65740 26628 65796 26630
rect 65820 26628 65876 26630
rect 65900 26628 65956 26630
rect 65660 25594 65716 25596
rect 65740 25594 65796 25596
rect 65820 25594 65876 25596
rect 65900 25594 65956 25596
rect 65660 25542 65706 25594
rect 65706 25542 65716 25594
rect 65740 25542 65770 25594
rect 65770 25542 65782 25594
rect 65782 25542 65796 25594
rect 65820 25542 65834 25594
rect 65834 25542 65846 25594
rect 65846 25542 65876 25594
rect 65900 25542 65910 25594
rect 65910 25542 65956 25594
rect 65660 25540 65716 25542
rect 65740 25540 65796 25542
rect 65820 25540 65876 25542
rect 65900 25540 65956 25542
rect 65660 24506 65716 24508
rect 65740 24506 65796 24508
rect 65820 24506 65876 24508
rect 65900 24506 65956 24508
rect 65660 24454 65706 24506
rect 65706 24454 65716 24506
rect 65740 24454 65770 24506
rect 65770 24454 65782 24506
rect 65782 24454 65796 24506
rect 65820 24454 65834 24506
rect 65834 24454 65846 24506
rect 65846 24454 65876 24506
rect 65900 24454 65910 24506
rect 65910 24454 65956 24506
rect 65660 24452 65716 24454
rect 65740 24452 65796 24454
rect 65820 24452 65876 24454
rect 65900 24452 65956 24454
rect 65660 23418 65716 23420
rect 65740 23418 65796 23420
rect 65820 23418 65876 23420
rect 65900 23418 65956 23420
rect 65660 23366 65706 23418
rect 65706 23366 65716 23418
rect 65740 23366 65770 23418
rect 65770 23366 65782 23418
rect 65782 23366 65796 23418
rect 65820 23366 65834 23418
rect 65834 23366 65846 23418
rect 65846 23366 65876 23418
rect 65900 23366 65910 23418
rect 65910 23366 65956 23418
rect 65660 23364 65716 23366
rect 65740 23364 65796 23366
rect 65820 23364 65876 23366
rect 65900 23364 65956 23366
rect 65660 22330 65716 22332
rect 65740 22330 65796 22332
rect 65820 22330 65876 22332
rect 65900 22330 65956 22332
rect 65660 22278 65706 22330
rect 65706 22278 65716 22330
rect 65740 22278 65770 22330
rect 65770 22278 65782 22330
rect 65782 22278 65796 22330
rect 65820 22278 65834 22330
rect 65834 22278 65846 22330
rect 65846 22278 65876 22330
rect 65900 22278 65910 22330
rect 65910 22278 65956 22330
rect 65660 22276 65716 22278
rect 65740 22276 65796 22278
rect 65820 22276 65876 22278
rect 65900 22276 65956 22278
rect 65660 21242 65716 21244
rect 65740 21242 65796 21244
rect 65820 21242 65876 21244
rect 65900 21242 65956 21244
rect 65660 21190 65706 21242
rect 65706 21190 65716 21242
rect 65740 21190 65770 21242
rect 65770 21190 65782 21242
rect 65782 21190 65796 21242
rect 65820 21190 65834 21242
rect 65834 21190 65846 21242
rect 65846 21190 65876 21242
rect 65900 21190 65910 21242
rect 65910 21190 65956 21242
rect 65660 21188 65716 21190
rect 65740 21188 65796 21190
rect 65820 21188 65876 21190
rect 65900 21188 65956 21190
rect 65660 20154 65716 20156
rect 65740 20154 65796 20156
rect 65820 20154 65876 20156
rect 65900 20154 65956 20156
rect 65660 20102 65706 20154
rect 65706 20102 65716 20154
rect 65740 20102 65770 20154
rect 65770 20102 65782 20154
rect 65782 20102 65796 20154
rect 65820 20102 65834 20154
rect 65834 20102 65846 20154
rect 65846 20102 65876 20154
rect 65900 20102 65910 20154
rect 65910 20102 65956 20154
rect 65660 20100 65716 20102
rect 65740 20100 65796 20102
rect 65820 20100 65876 20102
rect 65900 20100 65956 20102
rect 65660 19066 65716 19068
rect 65740 19066 65796 19068
rect 65820 19066 65876 19068
rect 65900 19066 65956 19068
rect 65660 19014 65706 19066
rect 65706 19014 65716 19066
rect 65740 19014 65770 19066
rect 65770 19014 65782 19066
rect 65782 19014 65796 19066
rect 65820 19014 65834 19066
rect 65834 19014 65846 19066
rect 65846 19014 65876 19066
rect 65900 19014 65910 19066
rect 65910 19014 65956 19066
rect 65660 19012 65716 19014
rect 65740 19012 65796 19014
rect 65820 19012 65876 19014
rect 65900 19012 65956 19014
rect 65660 17978 65716 17980
rect 65740 17978 65796 17980
rect 65820 17978 65876 17980
rect 65900 17978 65956 17980
rect 65660 17926 65706 17978
rect 65706 17926 65716 17978
rect 65740 17926 65770 17978
rect 65770 17926 65782 17978
rect 65782 17926 65796 17978
rect 65820 17926 65834 17978
rect 65834 17926 65846 17978
rect 65846 17926 65876 17978
rect 65900 17926 65910 17978
rect 65910 17926 65956 17978
rect 65660 17924 65716 17926
rect 65740 17924 65796 17926
rect 65820 17924 65876 17926
rect 65900 17924 65956 17926
rect 65660 16890 65716 16892
rect 65740 16890 65796 16892
rect 65820 16890 65876 16892
rect 65900 16890 65956 16892
rect 65660 16838 65706 16890
rect 65706 16838 65716 16890
rect 65740 16838 65770 16890
rect 65770 16838 65782 16890
rect 65782 16838 65796 16890
rect 65820 16838 65834 16890
rect 65834 16838 65846 16890
rect 65846 16838 65876 16890
rect 65900 16838 65910 16890
rect 65910 16838 65956 16890
rect 65660 16836 65716 16838
rect 65740 16836 65796 16838
rect 65820 16836 65876 16838
rect 65900 16836 65956 16838
rect 50300 16346 50356 16348
rect 50380 16346 50436 16348
rect 50460 16346 50516 16348
rect 50540 16346 50596 16348
rect 50300 16294 50346 16346
rect 50346 16294 50356 16346
rect 50380 16294 50410 16346
rect 50410 16294 50422 16346
rect 50422 16294 50436 16346
rect 50460 16294 50474 16346
rect 50474 16294 50486 16346
rect 50486 16294 50516 16346
rect 50540 16294 50550 16346
rect 50550 16294 50596 16346
rect 50300 16292 50356 16294
rect 50380 16292 50436 16294
rect 50460 16292 50516 16294
rect 50540 16292 50596 16294
rect 65660 15802 65716 15804
rect 65740 15802 65796 15804
rect 65820 15802 65876 15804
rect 65900 15802 65956 15804
rect 65660 15750 65706 15802
rect 65706 15750 65716 15802
rect 65740 15750 65770 15802
rect 65770 15750 65782 15802
rect 65782 15750 65796 15802
rect 65820 15750 65834 15802
rect 65834 15750 65846 15802
rect 65846 15750 65876 15802
rect 65900 15750 65910 15802
rect 65910 15750 65956 15802
rect 65660 15748 65716 15750
rect 65740 15748 65796 15750
rect 65820 15748 65876 15750
rect 65900 15748 65956 15750
rect 50300 15258 50356 15260
rect 50380 15258 50436 15260
rect 50460 15258 50516 15260
rect 50540 15258 50596 15260
rect 50300 15206 50346 15258
rect 50346 15206 50356 15258
rect 50380 15206 50410 15258
rect 50410 15206 50422 15258
rect 50422 15206 50436 15258
rect 50460 15206 50474 15258
rect 50474 15206 50486 15258
rect 50486 15206 50516 15258
rect 50540 15206 50550 15258
rect 50550 15206 50596 15258
rect 50300 15204 50356 15206
rect 50380 15204 50436 15206
rect 50460 15204 50516 15206
rect 50540 15204 50596 15206
rect 65660 14714 65716 14716
rect 65740 14714 65796 14716
rect 65820 14714 65876 14716
rect 65900 14714 65956 14716
rect 65660 14662 65706 14714
rect 65706 14662 65716 14714
rect 65740 14662 65770 14714
rect 65770 14662 65782 14714
rect 65782 14662 65796 14714
rect 65820 14662 65834 14714
rect 65834 14662 65846 14714
rect 65846 14662 65876 14714
rect 65900 14662 65910 14714
rect 65910 14662 65956 14714
rect 65660 14660 65716 14662
rect 65740 14660 65796 14662
rect 65820 14660 65876 14662
rect 65900 14660 65956 14662
rect 50300 14170 50356 14172
rect 50380 14170 50436 14172
rect 50460 14170 50516 14172
rect 50540 14170 50596 14172
rect 50300 14118 50346 14170
rect 50346 14118 50356 14170
rect 50380 14118 50410 14170
rect 50410 14118 50422 14170
rect 50422 14118 50436 14170
rect 50460 14118 50474 14170
rect 50474 14118 50486 14170
rect 50486 14118 50516 14170
rect 50540 14118 50550 14170
rect 50550 14118 50596 14170
rect 50300 14116 50356 14118
rect 50380 14116 50436 14118
rect 50460 14116 50516 14118
rect 50540 14116 50596 14118
rect 65660 13626 65716 13628
rect 65740 13626 65796 13628
rect 65820 13626 65876 13628
rect 65900 13626 65956 13628
rect 65660 13574 65706 13626
rect 65706 13574 65716 13626
rect 65740 13574 65770 13626
rect 65770 13574 65782 13626
rect 65782 13574 65796 13626
rect 65820 13574 65834 13626
rect 65834 13574 65846 13626
rect 65846 13574 65876 13626
rect 65900 13574 65910 13626
rect 65910 13574 65956 13626
rect 65660 13572 65716 13574
rect 65740 13572 65796 13574
rect 65820 13572 65876 13574
rect 65900 13572 65956 13574
rect 50300 13082 50356 13084
rect 50380 13082 50436 13084
rect 50460 13082 50516 13084
rect 50540 13082 50596 13084
rect 50300 13030 50346 13082
rect 50346 13030 50356 13082
rect 50380 13030 50410 13082
rect 50410 13030 50422 13082
rect 50422 13030 50436 13082
rect 50460 13030 50474 13082
rect 50474 13030 50486 13082
rect 50486 13030 50516 13082
rect 50540 13030 50550 13082
rect 50550 13030 50596 13082
rect 50300 13028 50356 13030
rect 50380 13028 50436 13030
rect 50460 13028 50516 13030
rect 50540 13028 50596 13030
rect 65660 12538 65716 12540
rect 65740 12538 65796 12540
rect 65820 12538 65876 12540
rect 65900 12538 65956 12540
rect 65660 12486 65706 12538
rect 65706 12486 65716 12538
rect 65740 12486 65770 12538
rect 65770 12486 65782 12538
rect 65782 12486 65796 12538
rect 65820 12486 65834 12538
rect 65834 12486 65846 12538
rect 65846 12486 65876 12538
rect 65900 12486 65910 12538
rect 65910 12486 65956 12538
rect 65660 12484 65716 12486
rect 65740 12484 65796 12486
rect 65820 12484 65876 12486
rect 65900 12484 65956 12486
rect 50300 11994 50356 11996
rect 50380 11994 50436 11996
rect 50460 11994 50516 11996
rect 50540 11994 50596 11996
rect 50300 11942 50346 11994
rect 50346 11942 50356 11994
rect 50380 11942 50410 11994
rect 50410 11942 50422 11994
rect 50422 11942 50436 11994
rect 50460 11942 50474 11994
rect 50474 11942 50486 11994
rect 50486 11942 50516 11994
rect 50540 11942 50550 11994
rect 50550 11942 50596 11994
rect 50300 11940 50356 11942
rect 50380 11940 50436 11942
rect 50460 11940 50516 11942
rect 50540 11940 50596 11942
rect 65660 11450 65716 11452
rect 65740 11450 65796 11452
rect 65820 11450 65876 11452
rect 65900 11450 65956 11452
rect 65660 11398 65706 11450
rect 65706 11398 65716 11450
rect 65740 11398 65770 11450
rect 65770 11398 65782 11450
rect 65782 11398 65796 11450
rect 65820 11398 65834 11450
rect 65834 11398 65846 11450
rect 65846 11398 65876 11450
rect 65900 11398 65910 11450
rect 65910 11398 65956 11450
rect 65660 11396 65716 11398
rect 65740 11396 65796 11398
rect 65820 11396 65876 11398
rect 65900 11396 65956 11398
rect 50300 10906 50356 10908
rect 50380 10906 50436 10908
rect 50460 10906 50516 10908
rect 50540 10906 50596 10908
rect 50300 10854 50346 10906
rect 50346 10854 50356 10906
rect 50380 10854 50410 10906
rect 50410 10854 50422 10906
rect 50422 10854 50436 10906
rect 50460 10854 50474 10906
rect 50474 10854 50486 10906
rect 50486 10854 50516 10906
rect 50540 10854 50550 10906
rect 50550 10854 50596 10906
rect 50300 10852 50356 10854
rect 50380 10852 50436 10854
rect 50460 10852 50516 10854
rect 50540 10852 50596 10854
rect 65660 10362 65716 10364
rect 65740 10362 65796 10364
rect 65820 10362 65876 10364
rect 65900 10362 65956 10364
rect 65660 10310 65706 10362
rect 65706 10310 65716 10362
rect 65740 10310 65770 10362
rect 65770 10310 65782 10362
rect 65782 10310 65796 10362
rect 65820 10310 65834 10362
rect 65834 10310 65846 10362
rect 65846 10310 65876 10362
rect 65900 10310 65910 10362
rect 65910 10310 65956 10362
rect 65660 10308 65716 10310
rect 65740 10308 65796 10310
rect 65820 10308 65876 10310
rect 65900 10308 65956 10310
rect 50300 9818 50356 9820
rect 50380 9818 50436 9820
rect 50460 9818 50516 9820
rect 50540 9818 50596 9820
rect 50300 9766 50346 9818
rect 50346 9766 50356 9818
rect 50380 9766 50410 9818
rect 50410 9766 50422 9818
rect 50422 9766 50436 9818
rect 50460 9766 50474 9818
rect 50474 9766 50486 9818
rect 50486 9766 50516 9818
rect 50540 9766 50550 9818
rect 50550 9766 50596 9818
rect 50300 9764 50356 9766
rect 50380 9764 50436 9766
rect 50460 9764 50516 9766
rect 50540 9764 50596 9766
rect 65660 9274 65716 9276
rect 65740 9274 65796 9276
rect 65820 9274 65876 9276
rect 65900 9274 65956 9276
rect 65660 9222 65706 9274
rect 65706 9222 65716 9274
rect 65740 9222 65770 9274
rect 65770 9222 65782 9274
rect 65782 9222 65796 9274
rect 65820 9222 65834 9274
rect 65834 9222 65846 9274
rect 65846 9222 65876 9274
rect 65900 9222 65910 9274
rect 65910 9222 65956 9274
rect 65660 9220 65716 9222
rect 65740 9220 65796 9222
rect 65820 9220 65876 9222
rect 65900 9220 65956 9222
rect 50300 8730 50356 8732
rect 50380 8730 50436 8732
rect 50460 8730 50516 8732
rect 50540 8730 50596 8732
rect 50300 8678 50346 8730
rect 50346 8678 50356 8730
rect 50380 8678 50410 8730
rect 50410 8678 50422 8730
rect 50422 8678 50436 8730
rect 50460 8678 50474 8730
rect 50474 8678 50486 8730
rect 50486 8678 50516 8730
rect 50540 8678 50550 8730
rect 50550 8678 50596 8730
rect 50300 8676 50356 8678
rect 50380 8676 50436 8678
rect 50460 8676 50516 8678
rect 50540 8676 50596 8678
rect 65660 8186 65716 8188
rect 65740 8186 65796 8188
rect 65820 8186 65876 8188
rect 65900 8186 65956 8188
rect 65660 8134 65706 8186
rect 65706 8134 65716 8186
rect 65740 8134 65770 8186
rect 65770 8134 65782 8186
rect 65782 8134 65796 8186
rect 65820 8134 65834 8186
rect 65834 8134 65846 8186
rect 65846 8134 65876 8186
rect 65900 8134 65910 8186
rect 65910 8134 65956 8186
rect 65660 8132 65716 8134
rect 65740 8132 65796 8134
rect 65820 8132 65876 8134
rect 65900 8132 65956 8134
rect 50300 7642 50356 7644
rect 50380 7642 50436 7644
rect 50460 7642 50516 7644
rect 50540 7642 50596 7644
rect 50300 7590 50346 7642
rect 50346 7590 50356 7642
rect 50380 7590 50410 7642
rect 50410 7590 50422 7642
rect 50422 7590 50436 7642
rect 50460 7590 50474 7642
rect 50474 7590 50486 7642
rect 50486 7590 50516 7642
rect 50540 7590 50550 7642
rect 50550 7590 50596 7642
rect 50300 7588 50356 7590
rect 50380 7588 50436 7590
rect 50460 7588 50516 7590
rect 50540 7588 50596 7590
rect 65660 7098 65716 7100
rect 65740 7098 65796 7100
rect 65820 7098 65876 7100
rect 65900 7098 65956 7100
rect 65660 7046 65706 7098
rect 65706 7046 65716 7098
rect 65740 7046 65770 7098
rect 65770 7046 65782 7098
rect 65782 7046 65796 7098
rect 65820 7046 65834 7098
rect 65834 7046 65846 7098
rect 65846 7046 65876 7098
rect 65900 7046 65910 7098
rect 65910 7046 65956 7098
rect 65660 7044 65716 7046
rect 65740 7044 65796 7046
rect 65820 7044 65876 7046
rect 65900 7044 65956 7046
rect 50300 6554 50356 6556
rect 50380 6554 50436 6556
rect 50460 6554 50516 6556
rect 50540 6554 50596 6556
rect 50300 6502 50346 6554
rect 50346 6502 50356 6554
rect 50380 6502 50410 6554
rect 50410 6502 50422 6554
rect 50422 6502 50436 6554
rect 50460 6502 50474 6554
rect 50474 6502 50486 6554
rect 50486 6502 50516 6554
rect 50540 6502 50550 6554
rect 50550 6502 50596 6554
rect 50300 6500 50356 6502
rect 50380 6500 50436 6502
rect 50460 6500 50516 6502
rect 50540 6500 50596 6502
rect 65660 6010 65716 6012
rect 65740 6010 65796 6012
rect 65820 6010 65876 6012
rect 65900 6010 65956 6012
rect 65660 5958 65706 6010
rect 65706 5958 65716 6010
rect 65740 5958 65770 6010
rect 65770 5958 65782 6010
rect 65782 5958 65796 6010
rect 65820 5958 65834 6010
rect 65834 5958 65846 6010
rect 65846 5958 65876 6010
rect 65900 5958 65910 6010
rect 65910 5958 65956 6010
rect 65660 5956 65716 5958
rect 65740 5956 65796 5958
rect 65820 5956 65876 5958
rect 65900 5956 65956 5958
rect 50300 5466 50356 5468
rect 50380 5466 50436 5468
rect 50460 5466 50516 5468
rect 50540 5466 50596 5468
rect 50300 5414 50346 5466
rect 50346 5414 50356 5466
rect 50380 5414 50410 5466
rect 50410 5414 50422 5466
rect 50422 5414 50436 5466
rect 50460 5414 50474 5466
rect 50474 5414 50486 5466
rect 50486 5414 50516 5466
rect 50540 5414 50550 5466
rect 50550 5414 50596 5466
rect 50300 5412 50356 5414
rect 50380 5412 50436 5414
rect 50460 5412 50516 5414
rect 50540 5412 50596 5414
rect 65660 4922 65716 4924
rect 65740 4922 65796 4924
rect 65820 4922 65876 4924
rect 65900 4922 65956 4924
rect 65660 4870 65706 4922
rect 65706 4870 65716 4922
rect 65740 4870 65770 4922
rect 65770 4870 65782 4922
rect 65782 4870 65796 4922
rect 65820 4870 65834 4922
rect 65834 4870 65846 4922
rect 65846 4870 65876 4922
rect 65900 4870 65910 4922
rect 65910 4870 65956 4922
rect 65660 4868 65716 4870
rect 65740 4868 65796 4870
rect 65820 4868 65876 4870
rect 65900 4868 65956 4870
rect 50300 4378 50356 4380
rect 50380 4378 50436 4380
rect 50460 4378 50516 4380
rect 50540 4378 50596 4380
rect 50300 4326 50346 4378
rect 50346 4326 50356 4378
rect 50380 4326 50410 4378
rect 50410 4326 50422 4378
rect 50422 4326 50436 4378
rect 50460 4326 50474 4378
rect 50474 4326 50486 4378
rect 50486 4326 50516 4378
rect 50540 4326 50550 4378
rect 50550 4326 50596 4378
rect 50300 4324 50356 4326
rect 50380 4324 50436 4326
rect 50460 4324 50516 4326
rect 50540 4324 50596 4326
rect 65660 3834 65716 3836
rect 65740 3834 65796 3836
rect 65820 3834 65876 3836
rect 65900 3834 65956 3836
rect 65660 3782 65706 3834
rect 65706 3782 65716 3834
rect 65740 3782 65770 3834
rect 65770 3782 65782 3834
rect 65782 3782 65796 3834
rect 65820 3782 65834 3834
rect 65834 3782 65846 3834
rect 65846 3782 65876 3834
rect 65900 3782 65910 3834
rect 65910 3782 65956 3834
rect 65660 3780 65716 3782
rect 65740 3780 65796 3782
rect 65820 3780 65876 3782
rect 65900 3780 65956 3782
rect 50300 3290 50356 3292
rect 50380 3290 50436 3292
rect 50460 3290 50516 3292
rect 50540 3290 50596 3292
rect 50300 3238 50346 3290
rect 50346 3238 50356 3290
rect 50380 3238 50410 3290
rect 50410 3238 50422 3290
rect 50422 3238 50436 3290
rect 50460 3238 50474 3290
rect 50474 3238 50486 3290
rect 50486 3238 50516 3290
rect 50540 3238 50550 3290
rect 50550 3238 50596 3290
rect 50300 3236 50356 3238
rect 50380 3236 50436 3238
rect 50460 3236 50516 3238
rect 50540 3236 50596 3238
rect 50300 2202 50356 2204
rect 50380 2202 50436 2204
rect 50460 2202 50516 2204
rect 50540 2202 50596 2204
rect 50300 2150 50346 2202
rect 50346 2150 50356 2202
rect 50380 2150 50410 2202
rect 50410 2150 50422 2202
rect 50422 2150 50436 2202
rect 50460 2150 50474 2202
rect 50474 2150 50486 2202
rect 50486 2150 50516 2202
rect 50540 2150 50550 2202
rect 50550 2150 50596 2202
rect 50300 2148 50356 2150
rect 50380 2148 50436 2150
rect 50460 2148 50516 2150
rect 50540 2148 50596 2150
rect 65660 2746 65716 2748
rect 65740 2746 65796 2748
rect 65820 2746 65876 2748
rect 65900 2746 65956 2748
rect 65660 2694 65706 2746
rect 65706 2694 65716 2746
rect 65740 2694 65770 2746
rect 65770 2694 65782 2746
rect 65782 2694 65796 2746
rect 65820 2694 65834 2746
rect 65834 2694 65846 2746
rect 65846 2694 65876 2746
rect 65900 2694 65910 2746
rect 65910 2694 65956 2746
rect 65660 2692 65716 2694
rect 65740 2692 65796 2694
rect 65820 2692 65876 2694
rect 65900 2692 65956 2694
rect 77206 12280 77262 12336
rect 77850 110200 77906 110256
rect 77850 106156 77852 106176
rect 77852 106156 77904 106176
rect 77904 106156 77906 106176
rect 77850 106120 77906 106156
rect 77850 102720 77906 102776
rect 77850 98660 77906 98696
rect 77850 98640 77852 98660
rect 77852 98640 77904 98660
rect 77904 98640 77906 98660
rect 78034 94560 78090 94616
rect 77942 90500 77998 90536
rect 77942 90480 77944 90500
rect 77944 90480 77996 90500
rect 77996 90480 77998 90500
rect 77942 87080 77998 87136
rect 77850 83000 77906 83056
rect 77850 71460 77906 71496
rect 77850 71440 77852 71460
rect 77852 71440 77904 71460
rect 77904 71440 77906 71460
rect 78034 74840 78090 74896
rect 77942 67360 77998 67416
rect 78034 63280 78090 63336
rect 77942 59200 77998 59256
rect 77850 55800 77906 55856
rect 77850 51756 77852 51776
rect 77852 51756 77904 51776
rect 77904 51756 77906 51776
rect 77850 51720 77906 51756
rect 78034 43596 78036 43616
rect 78036 43596 78088 43616
rect 78088 43596 78090 43616
rect 78034 43560 78090 43596
rect 78034 40160 78090 40216
rect 78034 36080 78090 36136
rect 77758 32000 77814 32056
rect 77942 27920 77998 27976
rect 77850 24556 77852 24576
rect 77852 24556 77904 24576
rect 77904 24556 77906 24576
rect 77850 24520 77906 24556
rect 78034 20440 78090 20496
rect 78034 16396 78036 16416
rect 78036 16396 78088 16416
rect 78088 16396 78090 16416
rect 78034 16360 78090 16396
rect 78034 8880 78090 8936
rect 77850 4800 77906 4856
rect 77666 720 77722 776
<< metal3 >>
rect 77201 118418 77267 118421
rect 79200 118418 80000 118448
rect 77201 118416 80000 118418
rect 77201 118360 77206 118416
rect 77262 118360 80000 118416
rect 77201 118358 80000 118360
rect 77201 118355 77267 118358
rect 79200 118328 80000 118358
rect 19568 117536 19888 117537
rect 19568 117472 19576 117536
rect 19640 117472 19656 117536
rect 19720 117472 19736 117536
rect 19800 117472 19816 117536
rect 19880 117472 19888 117536
rect 19568 117471 19888 117472
rect 50288 117536 50608 117537
rect 50288 117472 50296 117536
rect 50360 117472 50376 117536
rect 50440 117472 50456 117536
rect 50520 117472 50536 117536
rect 50600 117472 50608 117536
rect 50288 117471 50608 117472
rect 0 117058 800 117088
rect 1853 117058 1919 117061
rect 0 117056 1919 117058
rect 0 117000 1858 117056
rect 1914 117000 1919 117056
rect 0 116998 1919 117000
rect 0 116968 800 116998
rect 1853 116995 1919 116998
rect 4208 116992 4528 116993
rect 4208 116928 4216 116992
rect 4280 116928 4296 116992
rect 4360 116928 4376 116992
rect 4440 116928 4456 116992
rect 4520 116928 4528 116992
rect 4208 116927 4528 116928
rect 34928 116992 35248 116993
rect 34928 116928 34936 116992
rect 35000 116928 35016 116992
rect 35080 116928 35096 116992
rect 35160 116928 35176 116992
rect 35240 116928 35248 116992
rect 34928 116927 35248 116928
rect 65648 116992 65968 116993
rect 65648 116928 65656 116992
rect 65720 116928 65736 116992
rect 65800 116928 65816 116992
rect 65880 116928 65896 116992
rect 65960 116928 65968 116992
rect 65648 116927 65968 116928
rect 19568 116448 19888 116449
rect 19568 116384 19576 116448
rect 19640 116384 19656 116448
rect 19720 116384 19736 116448
rect 19800 116384 19816 116448
rect 19880 116384 19888 116448
rect 19568 116383 19888 116384
rect 50288 116448 50608 116449
rect 50288 116384 50296 116448
rect 50360 116384 50376 116448
rect 50440 116384 50456 116448
rect 50520 116384 50536 116448
rect 50600 116384 50608 116448
rect 50288 116383 50608 116384
rect 4208 115904 4528 115905
rect 4208 115840 4216 115904
rect 4280 115840 4296 115904
rect 4360 115840 4376 115904
rect 4440 115840 4456 115904
rect 4520 115840 4528 115904
rect 4208 115839 4528 115840
rect 34928 115904 35248 115905
rect 34928 115840 34936 115904
rect 35000 115840 35016 115904
rect 35080 115840 35096 115904
rect 35160 115840 35176 115904
rect 35240 115840 35248 115904
rect 34928 115839 35248 115840
rect 65648 115904 65968 115905
rect 65648 115840 65656 115904
rect 65720 115840 65736 115904
rect 65800 115840 65816 115904
rect 65880 115840 65896 115904
rect 65960 115840 65968 115904
rect 65648 115839 65968 115840
rect 19568 115360 19888 115361
rect 19568 115296 19576 115360
rect 19640 115296 19656 115360
rect 19720 115296 19736 115360
rect 19800 115296 19816 115360
rect 19880 115296 19888 115360
rect 19568 115295 19888 115296
rect 50288 115360 50608 115361
rect 50288 115296 50296 115360
rect 50360 115296 50376 115360
rect 50440 115296 50456 115360
rect 50520 115296 50536 115360
rect 50600 115296 50608 115360
rect 50288 115295 50608 115296
rect 4208 114816 4528 114817
rect 4208 114752 4216 114816
rect 4280 114752 4296 114816
rect 4360 114752 4376 114816
rect 4440 114752 4456 114816
rect 4520 114752 4528 114816
rect 4208 114751 4528 114752
rect 34928 114816 35248 114817
rect 34928 114752 34936 114816
rect 35000 114752 35016 114816
rect 35080 114752 35096 114816
rect 35160 114752 35176 114816
rect 35240 114752 35248 114816
rect 34928 114751 35248 114752
rect 65648 114816 65968 114817
rect 65648 114752 65656 114816
rect 65720 114752 65736 114816
rect 65800 114752 65816 114816
rect 65880 114752 65896 114816
rect 65960 114752 65968 114816
rect 65648 114751 65968 114752
rect 78029 114338 78095 114341
rect 79200 114338 80000 114368
rect 78029 114336 80000 114338
rect 78029 114280 78034 114336
rect 78090 114280 80000 114336
rect 78029 114278 80000 114280
rect 78029 114275 78095 114278
rect 19568 114272 19888 114273
rect 19568 114208 19576 114272
rect 19640 114208 19656 114272
rect 19720 114208 19736 114272
rect 19800 114208 19816 114272
rect 19880 114208 19888 114272
rect 19568 114207 19888 114208
rect 50288 114272 50608 114273
rect 50288 114208 50296 114272
rect 50360 114208 50376 114272
rect 50440 114208 50456 114272
rect 50520 114208 50536 114272
rect 50600 114208 50608 114272
rect 79200 114248 80000 114278
rect 50288 114207 50608 114208
rect 4208 113728 4528 113729
rect 4208 113664 4216 113728
rect 4280 113664 4296 113728
rect 4360 113664 4376 113728
rect 4440 113664 4456 113728
rect 4520 113664 4528 113728
rect 4208 113663 4528 113664
rect 34928 113728 35248 113729
rect 34928 113664 34936 113728
rect 35000 113664 35016 113728
rect 35080 113664 35096 113728
rect 35160 113664 35176 113728
rect 35240 113664 35248 113728
rect 34928 113663 35248 113664
rect 65648 113728 65968 113729
rect 65648 113664 65656 113728
rect 65720 113664 65736 113728
rect 65800 113664 65816 113728
rect 65880 113664 65896 113728
rect 65960 113664 65968 113728
rect 65648 113663 65968 113664
rect 19568 113184 19888 113185
rect 19568 113120 19576 113184
rect 19640 113120 19656 113184
rect 19720 113120 19736 113184
rect 19800 113120 19816 113184
rect 19880 113120 19888 113184
rect 19568 113119 19888 113120
rect 50288 113184 50608 113185
rect 50288 113120 50296 113184
rect 50360 113120 50376 113184
rect 50440 113120 50456 113184
rect 50520 113120 50536 113184
rect 50600 113120 50608 113184
rect 50288 113119 50608 113120
rect 0 112978 800 113008
rect 1577 112978 1643 112981
rect 0 112976 1643 112978
rect 0 112920 1582 112976
rect 1638 112920 1643 112976
rect 0 112918 1643 112920
rect 0 112888 800 112918
rect 1577 112915 1643 112918
rect 4208 112640 4528 112641
rect 4208 112576 4216 112640
rect 4280 112576 4296 112640
rect 4360 112576 4376 112640
rect 4440 112576 4456 112640
rect 4520 112576 4528 112640
rect 4208 112575 4528 112576
rect 34928 112640 35248 112641
rect 34928 112576 34936 112640
rect 35000 112576 35016 112640
rect 35080 112576 35096 112640
rect 35160 112576 35176 112640
rect 35240 112576 35248 112640
rect 34928 112575 35248 112576
rect 65648 112640 65968 112641
rect 65648 112576 65656 112640
rect 65720 112576 65736 112640
rect 65800 112576 65816 112640
rect 65880 112576 65896 112640
rect 65960 112576 65968 112640
rect 65648 112575 65968 112576
rect 19568 112096 19888 112097
rect 19568 112032 19576 112096
rect 19640 112032 19656 112096
rect 19720 112032 19736 112096
rect 19800 112032 19816 112096
rect 19880 112032 19888 112096
rect 19568 112031 19888 112032
rect 50288 112096 50608 112097
rect 50288 112032 50296 112096
rect 50360 112032 50376 112096
rect 50440 112032 50456 112096
rect 50520 112032 50536 112096
rect 50600 112032 50608 112096
rect 50288 112031 50608 112032
rect 4208 111552 4528 111553
rect 4208 111488 4216 111552
rect 4280 111488 4296 111552
rect 4360 111488 4376 111552
rect 4440 111488 4456 111552
rect 4520 111488 4528 111552
rect 4208 111487 4528 111488
rect 34928 111552 35248 111553
rect 34928 111488 34936 111552
rect 35000 111488 35016 111552
rect 35080 111488 35096 111552
rect 35160 111488 35176 111552
rect 35240 111488 35248 111552
rect 34928 111487 35248 111488
rect 65648 111552 65968 111553
rect 65648 111488 65656 111552
rect 65720 111488 65736 111552
rect 65800 111488 65816 111552
rect 65880 111488 65896 111552
rect 65960 111488 65968 111552
rect 65648 111487 65968 111488
rect 19568 111008 19888 111009
rect 19568 110944 19576 111008
rect 19640 110944 19656 111008
rect 19720 110944 19736 111008
rect 19800 110944 19816 111008
rect 19880 110944 19888 111008
rect 19568 110943 19888 110944
rect 50288 111008 50608 111009
rect 50288 110944 50296 111008
rect 50360 110944 50376 111008
rect 50440 110944 50456 111008
rect 50520 110944 50536 111008
rect 50600 110944 50608 111008
rect 50288 110943 50608 110944
rect 4208 110464 4528 110465
rect 4208 110400 4216 110464
rect 4280 110400 4296 110464
rect 4360 110400 4376 110464
rect 4440 110400 4456 110464
rect 4520 110400 4528 110464
rect 4208 110399 4528 110400
rect 34928 110464 35248 110465
rect 34928 110400 34936 110464
rect 35000 110400 35016 110464
rect 35080 110400 35096 110464
rect 35160 110400 35176 110464
rect 35240 110400 35248 110464
rect 34928 110399 35248 110400
rect 65648 110464 65968 110465
rect 65648 110400 65656 110464
rect 65720 110400 65736 110464
rect 65800 110400 65816 110464
rect 65880 110400 65896 110464
rect 65960 110400 65968 110464
rect 65648 110399 65968 110400
rect 77845 110258 77911 110261
rect 79200 110258 80000 110288
rect 77845 110256 80000 110258
rect 77845 110200 77850 110256
rect 77906 110200 80000 110256
rect 77845 110198 80000 110200
rect 77845 110195 77911 110198
rect 79200 110168 80000 110198
rect 19568 109920 19888 109921
rect 19568 109856 19576 109920
rect 19640 109856 19656 109920
rect 19720 109856 19736 109920
rect 19800 109856 19816 109920
rect 19880 109856 19888 109920
rect 19568 109855 19888 109856
rect 50288 109920 50608 109921
rect 50288 109856 50296 109920
rect 50360 109856 50376 109920
rect 50440 109856 50456 109920
rect 50520 109856 50536 109920
rect 50600 109856 50608 109920
rect 50288 109855 50608 109856
rect 0 109578 800 109608
rect 1853 109578 1919 109581
rect 0 109576 1919 109578
rect 0 109520 1858 109576
rect 1914 109520 1919 109576
rect 0 109518 1919 109520
rect 0 109488 800 109518
rect 1853 109515 1919 109518
rect 4208 109376 4528 109377
rect 4208 109312 4216 109376
rect 4280 109312 4296 109376
rect 4360 109312 4376 109376
rect 4440 109312 4456 109376
rect 4520 109312 4528 109376
rect 4208 109311 4528 109312
rect 34928 109376 35248 109377
rect 34928 109312 34936 109376
rect 35000 109312 35016 109376
rect 35080 109312 35096 109376
rect 35160 109312 35176 109376
rect 35240 109312 35248 109376
rect 34928 109311 35248 109312
rect 65648 109376 65968 109377
rect 65648 109312 65656 109376
rect 65720 109312 65736 109376
rect 65800 109312 65816 109376
rect 65880 109312 65896 109376
rect 65960 109312 65968 109376
rect 65648 109311 65968 109312
rect 19568 108832 19888 108833
rect 19568 108768 19576 108832
rect 19640 108768 19656 108832
rect 19720 108768 19736 108832
rect 19800 108768 19816 108832
rect 19880 108768 19888 108832
rect 19568 108767 19888 108768
rect 50288 108832 50608 108833
rect 50288 108768 50296 108832
rect 50360 108768 50376 108832
rect 50440 108768 50456 108832
rect 50520 108768 50536 108832
rect 50600 108768 50608 108832
rect 50288 108767 50608 108768
rect 4208 108288 4528 108289
rect 4208 108224 4216 108288
rect 4280 108224 4296 108288
rect 4360 108224 4376 108288
rect 4440 108224 4456 108288
rect 4520 108224 4528 108288
rect 4208 108223 4528 108224
rect 34928 108288 35248 108289
rect 34928 108224 34936 108288
rect 35000 108224 35016 108288
rect 35080 108224 35096 108288
rect 35160 108224 35176 108288
rect 35240 108224 35248 108288
rect 34928 108223 35248 108224
rect 65648 108288 65968 108289
rect 65648 108224 65656 108288
rect 65720 108224 65736 108288
rect 65800 108224 65816 108288
rect 65880 108224 65896 108288
rect 65960 108224 65968 108288
rect 65648 108223 65968 108224
rect 19568 107744 19888 107745
rect 19568 107680 19576 107744
rect 19640 107680 19656 107744
rect 19720 107680 19736 107744
rect 19800 107680 19816 107744
rect 19880 107680 19888 107744
rect 19568 107679 19888 107680
rect 50288 107744 50608 107745
rect 50288 107680 50296 107744
rect 50360 107680 50376 107744
rect 50440 107680 50456 107744
rect 50520 107680 50536 107744
rect 50600 107680 50608 107744
rect 50288 107679 50608 107680
rect 4208 107200 4528 107201
rect 4208 107136 4216 107200
rect 4280 107136 4296 107200
rect 4360 107136 4376 107200
rect 4440 107136 4456 107200
rect 4520 107136 4528 107200
rect 4208 107135 4528 107136
rect 34928 107200 35248 107201
rect 34928 107136 34936 107200
rect 35000 107136 35016 107200
rect 35080 107136 35096 107200
rect 35160 107136 35176 107200
rect 35240 107136 35248 107200
rect 34928 107135 35248 107136
rect 65648 107200 65968 107201
rect 65648 107136 65656 107200
rect 65720 107136 65736 107200
rect 65800 107136 65816 107200
rect 65880 107136 65896 107200
rect 65960 107136 65968 107200
rect 65648 107135 65968 107136
rect 19568 106656 19888 106657
rect 19568 106592 19576 106656
rect 19640 106592 19656 106656
rect 19720 106592 19736 106656
rect 19800 106592 19816 106656
rect 19880 106592 19888 106656
rect 19568 106591 19888 106592
rect 50288 106656 50608 106657
rect 50288 106592 50296 106656
rect 50360 106592 50376 106656
rect 50440 106592 50456 106656
rect 50520 106592 50536 106656
rect 50600 106592 50608 106656
rect 50288 106591 50608 106592
rect 77845 106178 77911 106181
rect 79200 106178 80000 106208
rect 77845 106176 80000 106178
rect 77845 106120 77850 106176
rect 77906 106120 80000 106176
rect 77845 106118 80000 106120
rect 77845 106115 77911 106118
rect 4208 106112 4528 106113
rect 4208 106048 4216 106112
rect 4280 106048 4296 106112
rect 4360 106048 4376 106112
rect 4440 106048 4456 106112
rect 4520 106048 4528 106112
rect 4208 106047 4528 106048
rect 34928 106112 35248 106113
rect 34928 106048 34936 106112
rect 35000 106048 35016 106112
rect 35080 106048 35096 106112
rect 35160 106048 35176 106112
rect 35240 106048 35248 106112
rect 34928 106047 35248 106048
rect 65648 106112 65968 106113
rect 65648 106048 65656 106112
rect 65720 106048 65736 106112
rect 65800 106048 65816 106112
rect 65880 106048 65896 106112
rect 65960 106048 65968 106112
rect 79200 106088 80000 106118
rect 65648 106047 65968 106048
rect 19568 105568 19888 105569
rect 0 105498 800 105528
rect 19568 105504 19576 105568
rect 19640 105504 19656 105568
rect 19720 105504 19736 105568
rect 19800 105504 19816 105568
rect 19880 105504 19888 105568
rect 19568 105503 19888 105504
rect 50288 105568 50608 105569
rect 50288 105504 50296 105568
rect 50360 105504 50376 105568
rect 50440 105504 50456 105568
rect 50520 105504 50536 105568
rect 50600 105504 50608 105568
rect 50288 105503 50608 105504
rect 1393 105498 1459 105501
rect 0 105496 1459 105498
rect 0 105440 1398 105496
rect 1454 105440 1459 105496
rect 0 105438 1459 105440
rect 0 105408 800 105438
rect 1393 105435 1459 105438
rect 4208 105024 4528 105025
rect 4208 104960 4216 105024
rect 4280 104960 4296 105024
rect 4360 104960 4376 105024
rect 4440 104960 4456 105024
rect 4520 104960 4528 105024
rect 4208 104959 4528 104960
rect 34928 105024 35248 105025
rect 34928 104960 34936 105024
rect 35000 104960 35016 105024
rect 35080 104960 35096 105024
rect 35160 104960 35176 105024
rect 35240 104960 35248 105024
rect 34928 104959 35248 104960
rect 65648 105024 65968 105025
rect 65648 104960 65656 105024
rect 65720 104960 65736 105024
rect 65800 104960 65816 105024
rect 65880 104960 65896 105024
rect 65960 104960 65968 105024
rect 65648 104959 65968 104960
rect 19568 104480 19888 104481
rect 19568 104416 19576 104480
rect 19640 104416 19656 104480
rect 19720 104416 19736 104480
rect 19800 104416 19816 104480
rect 19880 104416 19888 104480
rect 19568 104415 19888 104416
rect 50288 104480 50608 104481
rect 50288 104416 50296 104480
rect 50360 104416 50376 104480
rect 50440 104416 50456 104480
rect 50520 104416 50536 104480
rect 50600 104416 50608 104480
rect 50288 104415 50608 104416
rect 4208 103936 4528 103937
rect 4208 103872 4216 103936
rect 4280 103872 4296 103936
rect 4360 103872 4376 103936
rect 4440 103872 4456 103936
rect 4520 103872 4528 103936
rect 4208 103871 4528 103872
rect 34928 103936 35248 103937
rect 34928 103872 34936 103936
rect 35000 103872 35016 103936
rect 35080 103872 35096 103936
rect 35160 103872 35176 103936
rect 35240 103872 35248 103936
rect 34928 103871 35248 103872
rect 65648 103936 65968 103937
rect 65648 103872 65656 103936
rect 65720 103872 65736 103936
rect 65800 103872 65816 103936
rect 65880 103872 65896 103936
rect 65960 103872 65968 103936
rect 65648 103871 65968 103872
rect 19568 103392 19888 103393
rect 19568 103328 19576 103392
rect 19640 103328 19656 103392
rect 19720 103328 19736 103392
rect 19800 103328 19816 103392
rect 19880 103328 19888 103392
rect 19568 103327 19888 103328
rect 50288 103392 50608 103393
rect 50288 103328 50296 103392
rect 50360 103328 50376 103392
rect 50440 103328 50456 103392
rect 50520 103328 50536 103392
rect 50600 103328 50608 103392
rect 50288 103327 50608 103328
rect 4208 102848 4528 102849
rect 4208 102784 4216 102848
rect 4280 102784 4296 102848
rect 4360 102784 4376 102848
rect 4440 102784 4456 102848
rect 4520 102784 4528 102848
rect 4208 102783 4528 102784
rect 34928 102848 35248 102849
rect 34928 102784 34936 102848
rect 35000 102784 35016 102848
rect 35080 102784 35096 102848
rect 35160 102784 35176 102848
rect 35240 102784 35248 102848
rect 34928 102783 35248 102784
rect 65648 102848 65968 102849
rect 65648 102784 65656 102848
rect 65720 102784 65736 102848
rect 65800 102784 65816 102848
rect 65880 102784 65896 102848
rect 65960 102784 65968 102848
rect 65648 102783 65968 102784
rect 77845 102778 77911 102781
rect 79200 102778 80000 102808
rect 77845 102776 80000 102778
rect 77845 102720 77850 102776
rect 77906 102720 80000 102776
rect 77845 102718 80000 102720
rect 77845 102715 77911 102718
rect 79200 102688 80000 102718
rect 19568 102304 19888 102305
rect 19568 102240 19576 102304
rect 19640 102240 19656 102304
rect 19720 102240 19736 102304
rect 19800 102240 19816 102304
rect 19880 102240 19888 102304
rect 19568 102239 19888 102240
rect 50288 102304 50608 102305
rect 50288 102240 50296 102304
rect 50360 102240 50376 102304
rect 50440 102240 50456 102304
rect 50520 102240 50536 102304
rect 50600 102240 50608 102304
rect 50288 102239 50608 102240
rect 4208 101760 4528 101761
rect 4208 101696 4216 101760
rect 4280 101696 4296 101760
rect 4360 101696 4376 101760
rect 4440 101696 4456 101760
rect 4520 101696 4528 101760
rect 4208 101695 4528 101696
rect 34928 101760 35248 101761
rect 34928 101696 34936 101760
rect 35000 101696 35016 101760
rect 35080 101696 35096 101760
rect 35160 101696 35176 101760
rect 35240 101696 35248 101760
rect 34928 101695 35248 101696
rect 65648 101760 65968 101761
rect 65648 101696 65656 101760
rect 65720 101696 65736 101760
rect 65800 101696 65816 101760
rect 65880 101696 65896 101760
rect 65960 101696 65968 101760
rect 65648 101695 65968 101696
rect 0 101418 800 101448
rect 1393 101418 1459 101421
rect 0 101416 1459 101418
rect 0 101360 1398 101416
rect 1454 101360 1459 101416
rect 0 101358 1459 101360
rect 0 101328 800 101358
rect 1393 101355 1459 101358
rect 19568 101216 19888 101217
rect 19568 101152 19576 101216
rect 19640 101152 19656 101216
rect 19720 101152 19736 101216
rect 19800 101152 19816 101216
rect 19880 101152 19888 101216
rect 19568 101151 19888 101152
rect 50288 101216 50608 101217
rect 50288 101152 50296 101216
rect 50360 101152 50376 101216
rect 50440 101152 50456 101216
rect 50520 101152 50536 101216
rect 50600 101152 50608 101216
rect 50288 101151 50608 101152
rect 4208 100672 4528 100673
rect 4208 100608 4216 100672
rect 4280 100608 4296 100672
rect 4360 100608 4376 100672
rect 4440 100608 4456 100672
rect 4520 100608 4528 100672
rect 4208 100607 4528 100608
rect 34928 100672 35248 100673
rect 34928 100608 34936 100672
rect 35000 100608 35016 100672
rect 35080 100608 35096 100672
rect 35160 100608 35176 100672
rect 35240 100608 35248 100672
rect 34928 100607 35248 100608
rect 65648 100672 65968 100673
rect 65648 100608 65656 100672
rect 65720 100608 65736 100672
rect 65800 100608 65816 100672
rect 65880 100608 65896 100672
rect 65960 100608 65968 100672
rect 65648 100607 65968 100608
rect 19568 100128 19888 100129
rect 19568 100064 19576 100128
rect 19640 100064 19656 100128
rect 19720 100064 19736 100128
rect 19800 100064 19816 100128
rect 19880 100064 19888 100128
rect 19568 100063 19888 100064
rect 50288 100128 50608 100129
rect 50288 100064 50296 100128
rect 50360 100064 50376 100128
rect 50440 100064 50456 100128
rect 50520 100064 50536 100128
rect 50600 100064 50608 100128
rect 50288 100063 50608 100064
rect 4208 99584 4528 99585
rect 4208 99520 4216 99584
rect 4280 99520 4296 99584
rect 4360 99520 4376 99584
rect 4440 99520 4456 99584
rect 4520 99520 4528 99584
rect 4208 99519 4528 99520
rect 34928 99584 35248 99585
rect 34928 99520 34936 99584
rect 35000 99520 35016 99584
rect 35080 99520 35096 99584
rect 35160 99520 35176 99584
rect 35240 99520 35248 99584
rect 34928 99519 35248 99520
rect 65648 99584 65968 99585
rect 65648 99520 65656 99584
rect 65720 99520 65736 99584
rect 65800 99520 65816 99584
rect 65880 99520 65896 99584
rect 65960 99520 65968 99584
rect 65648 99519 65968 99520
rect 19568 99040 19888 99041
rect 19568 98976 19576 99040
rect 19640 98976 19656 99040
rect 19720 98976 19736 99040
rect 19800 98976 19816 99040
rect 19880 98976 19888 99040
rect 19568 98975 19888 98976
rect 50288 99040 50608 99041
rect 50288 98976 50296 99040
rect 50360 98976 50376 99040
rect 50440 98976 50456 99040
rect 50520 98976 50536 99040
rect 50600 98976 50608 99040
rect 50288 98975 50608 98976
rect 77845 98698 77911 98701
rect 79200 98698 80000 98728
rect 77845 98696 80000 98698
rect 77845 98640 77850 98696
rect 77906 98640 80000 98696
rect 77845 98638 80000 98640
rect 77845 98635 77911 98638
rect 79200 98608 80000 98638
rect 4208 98496 4528 98497
rect 4208 98432 4216 98496
rect 4280 98432 4296 98496
rect 4360 98432 4376 98496
rect 4440 98432 4456 98496
rect 4520 98432 4528 98496
rect 4208 98431 4528 98432
rect 34928 98496 35248 98497
rect 34928 98432 34936 98496
rect 35000 98432 35016 98496
rect 35080 98432 35096 98496
rect 35160 98432 35176 98496
rect 35240 98432 35248 98496
rect 34928 98431 35248 98432
rect 65648 98496 65968 98497
rect 65648 98432 65656 98496
rect 65720 98432 65736 98496
rect 65800 98432 65816 98496
rect 65880 98432 65896 98496
rect 65960 98432 65968 98496
rect 65648 98431 65968 98432
rect 19568 97952 19888 97953
rect 19568 97888 19576 97952
rect 19640 97888 19656 97952
rect 19720 97888 19736 97952
rect 19800 97888 19816 97952
rect 19880 97888 19888 97952
rect 19568 97887 19888 97888
rect 50288 97952 50608 97953
rect 50288 97888 50296 97952
rect 50360 97888 50376 97952
rect 50440 97888 50456 97952
rect 50520 97888 50536 97952
rect 50600 97888 50608 97952
rect 50288 97887 50608 97888
rect 4208 97408 4528 97409
rect 0 97338 800 97368
rect 4208 97344 4216 97408
rect 4280 97344 4296 97408
rect 4360 97344 4376 97408
rect 4440 97344 4456 97408
rect 4520 97344 4528 97408
rect 4208 97343 4528 97344
rect 34928 97408 35248 97409
rect 34928 97344 34936 97408
rect 35000 97344 35016 97408
rect 35080 97344 35096 97408
rect 35160 97344 35176 97408
rect 35240 97344 35248 97408
rect 34928 97343 35248 97344
rect 65648 97408 65968 97409
rect 65648 97344 65656 97408
rect 65720 97344 65736 97408
rect 65800 97344 65816 97408
rect 65880 97344 65896 97408
rect 65960 97344 65968 97408
rect 65648 97343 65968 97344
rect 1393 97338 1459 97341
rect 0 97336 1459 97338
rect 0 97280 1398 97336
rect 1454 97280 1459 97336
rect 0 97278 1459 97280
rect 0 97248 800 97278
rect 1393 97275 1459 97278
rect 19568 96864 19888 96865
rect 19568 96800 19576 96864
rect 19640 96800 19656 96864
rect 19720 96800 19736 96864
rect 19800 96800 19816 96864
rect 19880 96800 19888 96864
rect 19568 96799 19888 96800
rect 50288 96864 50608 96865
rect 50288 96800 50296 96864
rect 50360 96800 50376 96864
rect 50440 96800 50456 96864
rect 50520 96800 50536 96864
rect 50600 96800 50608 96864
rect 50288 96799 50608 96800
rect 4208 96320 4528 96321
rect 4208 96256 4216 96320
rect 4280 96256 4296 96320
rect 4360 96256 4376 96320
rect 4440 96256 4456 96320
rect 4520 96256 4528 96320
rect 4208 96255 4528 96256
rect 34928 96320 35248 96321
rect 34928 96256 34936 96320
rect 35000 96256 35016 96320
rect 35080 96256 35096 96320
rect 35160 96256 35176 96320
rect 35240 96256 35248 96320
rect 34928 96255 35248 96256
rect 65648 96320 65968 96321
rect 65648 96256 65656 96320
rect 65720 96256 65736 96320
rect 65800 96256 65816 96320
rect 65880 96256 65896 96320
rect 65960 96256 65968 96320
rect 65648 96255 65968 96256
rect 19568 95776 19888 95777
rect 19568 95712 19576 95776
rect 19640 95712 19656 95776
rect 19720 95712 19736 95776
rect 19800 95712 19816 95776
rect 19880 95712 19888 95776
rect 19568 95711 19888 95712
rect 50288 95776 50608 95777
rect 50288 95712 50296 95776
rect 50360 95712 50376 95776
rect 50440 95712 50456 95776
rect 50520 95712 50536 95776
rect 50600 95712 50608 95776
rect 50288 95711 50608 95712
rect 4208 95232 4528 95233
rect 4208 95168 4216 95232
rect 4280 95168 4296 95232
rect 4360 95168 4376 95232
rect 4440 95168 4456 95232
rect 4520 95168 4528 95232
rect 4208 95167 4528 95168
rect 34928 95232 35248 95233
rect 34928 95168 34936 95232
rect 35000 95168 35016 95232
rect 35080 95168 35096 95232
rect 35160 95168 35176 95232
rect 35240 95168 35248 95232
rect 34928 95167 35248 95168
rect 65648 95232 65968 95233
rect 65648 95168 65656 95232
rect 65720 95168 65736 95232
rect 65800 95168 65816 95232
rect 65880 95168 65896 95232
rect 65960 95168 65968 95232
rect 65648 95167 65968 95168
rect 19568 94688 19888 94689
rect 19568 94624 19576 94688
rect 19640 94624 19656 94688
rect 19720 94624 19736 94688
rect 19800 94624 19816 94688
rect 19880 94624 19888 94688
rect 19568 94623 19888 94624
rect 50288 94688 50608 94689
rect 50288 94624 50296 94688
rect 50360 94624 50376 94688
rect 50440 94624 50456 94688
rect 50520 94624 50536 94688
rect 50600 94624 50608 94688
rect 50288 94623 50608 94624
rect 78029 94618 78095 94621
rect 79200 94618 80000 94648
rect 78029 94616 80000 94618
rect 78029 94560 78034 94616
rect 78090 94560 80000 94616
rect 78029 94558 80000 94560
rect 78029 94555 78095 94558
rect 79200 94528 80000 94558
rect 4208 94144 4528 94145
rect 4208 94080 4216 94144
rect 4280 94080 4296 94144
rect 4360 94080 4376 94144
rect 4440 94080 4456 94144
rect 4520 94080 4528 94144
rect 4208 94079 4528 94080
rect 34928 94144 35248 94145
rect 34928 94080 34936 94144
rect 35000 94080 35016 94144
rect 35080 94080 35096 94144
rect 35160 94080 35176 94144
rect 35240 94080 35248 94144
rect 34928 94079 35248 94080
rect 65648 94144 65968 94145
rect 65648 94080 65656 94144
rect 65720 94080 65736 94144
rect 65800 94080 65816 94144
rect 65880 94080 65896 94144
rect 65960 94080 65968 94144
rect 65648 94079 65968 94080
rect 0 93938 800 93968
rect 1577 93938 1643 93941
rect 0 93936 1643 93938
rect 0 93880 1582 93936
rect 1638 93880 1643 93936
rect 0 93878 1643 93880
rect 0 93848 800 93878
rect 1577 93875 1643 93878
rect 19568 93600 19888 93601
rect 19568 93536 19576 93600
rect 19640 93536 19656 93600
rect 19720 93536 19736 93600
rect 19800 93536 19816 93600
rect 19880 93536 19888 93600
rect 19568 93535 19888 93536
rect 50288 93600 50608 93601
rect 50288 93536 50296 93600
rect 50360 93536 50376 93600
rect 50440 93536 50456 93600
rect 50520 93536 50536 93600
rect 50600 93536 50608 93600
rect 50288 93535 50608 93536
rect 4208 93056 4528 93057
rect 4208 92992 4216 93056
rect 4280 92992 4296 93056
rect 4360 92992 4376 93056
rect 4440 92992 4456 93056
rect 4520 92992 4528 93056
rect 4208 92991 4528 92992
rect 34928 93056 35248 93057
rect 34928 92992 34936 93056
rect 35000 92992 35016 93056
rect 35080 92992 35096 93056
rect 35160 92992 35176 93056
rect 35240 92992 35248 93056
rect 34928 92991 35248 92992
rect 65648 93056 65968 93057
rect 65648 92992 65656 93056
rect 65720 92992 65736 93056
rect 65800 92992 65816 93056
rect 65880 92992 65896 93056
rect 65960 92992 65968 93056
rect 65648 92991 65968 92992
rect 19568 92512 19888 92513
rect 19568 92448 19576 92512
rect 19640 92448 19656 92512
rect 19720 92448 19736 92512
rect 19800 92448 19816 92512
rect 19880 92448 19888 92512
rect 19568 92447 19888 92448
rect 50288 92512 50608 92513
rect 50288 92448 50296 92512
rect 50360 92448 50376 92512
rect 50440 92448 50456 92512
rect 50520 92448 50536 92512
rect 50600 92448 50608 92512
rect 50288 92447 50608 92448
rect 4208 91968 4528 91969
rect 4208 91904 4216 91968
rect 4280 91904 4296 91968
rect 4360 91904 4376 91968
rect 4440 91904 4456 91968
rect 4520 91904 4528 91968
rect 4208 91903 4528 91904
rect 34928 91968 35248 91969
rect 34928 91904 34936 91968
rect 35000 91904 35016 91968
rect 35080 91904 35096 91968
rect 35160 91904 35176 91968
rect 35240 91904 35248 91968
rect 34928 91903 35248 91904
rect 65648 91968 65968 91969
rect 65648 91904 65656 91968
rect 65720 91904 65736 91968
rect 65800 91904 65816 91968
rect 65880 91904 65896 91968
rect 65960 91904 65968 91968
rect 65648 91903 65968 91904
rect 19568 91424 19888 91425
rect 19568 91360 19576 91424
rect 19640 91360 19656 91424
rect 19720 91360 19736 91424
rect 19800 91360 19816 91424
rect 19880 91360 19888 91424
rect 19568 91359 19888 91360
rect 50288 91424 50608 91425
rect 50288 91360 50296 91424
rect 50360 91360 50376 91424
rect 50440 91360 50456 91424
rect 50520 91360 50536 91424
rect 50600 91360 50608 91424
rect 50288 91359 50608 91360
rect 4208 90880 4528 90881
rect 4208 90816 4216 90880
rect 4280 90816 4296 90880
rect 4360 90816 4376 90880
rect 4440 90816 4456 90880
rect 4520 90816 4528 90880
rect 4208 90815 4528 90816
rect 34928 90880 35248 90881
rect 34928 90816 34936 90880
rect 35000 90816 35016 90880
rect 35080 90816 35096 90880
rect 35160 90816 35176 90880
rect 35240 90816 35248 90880
rect 34928 90815 35248 90816
rect 65648 90880 65968 90881
rect 65648 90816 65656 90880
rect 65720 90816 65736 90880
rect 65800 90816 65816 90880
rect 65880 90816 65896 90880
rect 65960 90816 65968 90880
rect 65648 90815 65968 90816
rect 77937 90538 78003 90541
rect 79200 90538 80000 90568
rect 77937 90536 80000 90538
rect 77937 90480 77942 90536
rect 77998 90480 80000 90536
rect 77937 90478 80000 90480
rect 77937 90475 78003 90478
rect 79200 90448 80000 90478
rect 19568 90336 19888 90337
rect 19568 90272 19576 90336
rect 19640 90272 19656 90336
rect 19720 90272 19736 90336
rect 19800 90272 19816 90336
rect 19880 90272 19888 90336
rect 19568 90271 19888 90272
rect 50288 90336 50608 90337
rect 50288 90272 50296 90336
rect 50360 90272 50376 90336
rect 50440 90272 50456 90336
rect 50520 90272 50536 90336
rect 50600 90272 50608 90336
rect 50288 90271 50608 90272
rect 0 89858 800 89888
rect 1485 89858 1551 89861
rect 0 89856 1551 89858
rect 0 89800 1490 89856
rect 1546 89800 1551 89856
rect 0 89798 1551 89800
rect 0 89768 800 89798
rect 1485 89795 1551 89798
rect 4208 89792 4528 89793
rect 4208 89728 4216 89792
rect 4280 89728 4296 89792
rect 4360 89728 4376 89792
rect 4440 89728 4456 89792
rect 4520 89728 4528 89792
rect 4208 89727 4528 89728
rect 34928 89792 35248 89793
rect 34928 89728 34936 89792
rect 35000 89728 35016 89792
rect 35080 89728 35096 89792
rect 35160 89728 35176 89792
rect 35240 89728 35248 89792
rect 34928 89727 35248 89728
rect 65648 89792 65968 89793
rect 65648 89728 65656 89792
rect 65720 89728 65736 89792
rect 65800 89728 65816 89792
rect 65880 89728 65896 89792
rect 65960 89728 65968 89792
rect 65648 89727 65968 89728
rect 19568 89248 19888 89249
rect 19568 89184 19576 89248
rect 19640 89184 19656 89248
rect 19720 89184 19736 89248
rect 19800 89184 19816 89248
rect 19880 89184 19888 89248
rect 19568 89183 19888 89184
rect 50288 89248 50608 89249
rect 50288 89184 50296 89248
rect 50360 89184 50376 89248
rect 50440 89184 50456 89248
rect 50520 89184 50536 89248
rect 50600 89184 50608 89248
rect 50288 89183 50608 89184
rect 4208 88704 4528 88705
rect 4208 88640 4216 88704
rect 4280 88640 4296 88704
rect 4360 88640 4376 88704
rect 4440 88640 4456 88704
rect 4520 88640 4528 88704
rect 4208 88639 4528 88640
rect 34928 88704 35248 88705
rect 34928 88640 34936 88704
rect 35000 88640 35016 88704
rect 35080 88640 35096 88704
rect 35160 88640 35176 88704
rect 35240 88640 35248 88704
rect 34928 88639 35248 88640
rect 65648 88704 65968 88705
rect 65648 88640 65656 88704
rect 65720 88640 65736 88704
rect 65800 88640 65816 88704
rect 65880 88640 65896 88704
rect 65960 88640 65968 88704
rect 65648 88639 65968 88640
rect 19568 88160 19888 88161
rect 19568 88096 19576 88160
rect 19640 88096 19656 88160
rect 19720 88096 19736 88160
rect 19800 88096 19816 88160
rect 19880 88096 19888 88160
rect 19568 88095 19888 88096
rect 50288 88160 50608 88161
rect 50288 88096 50296 88160
rect 50360 88096 50376 88160
rect 50440 88096 50456 88160
rect 50520 88096 50536 88160
rect 50600 88096 50608 88160
rect 50288 88095 50608 88096
rect 4208 87616 4528 87617
rect 4208 87552 4216 87616
rect 4280 87552 4296 87616
rect 4360 87552 4376 87616
rect 4440 87552 4456 87616
rect 4520 87552 4528 87616
rect 4208 87551 4528 87552
rect 34928 87616 35248 87617
rect 34928 87552 34936 87616
rect 35000 87552 35016 87616
rect 35080 87552 35096 87616
rect 35160 87552 35176 87616
rect 35240 87552 35248 87616
rect 34928 87551 35248 87552
rect 65648 87616 65968 87617
rect 65648 87552 65656 87616
rect 65720 87552 65736 87616
rect 65800 87552 65816 87616
rect 65880 87552 65896 87616
rect 65960 87552 65968 87616
rect 65648 87551 65968 87552
rect 77937 87138 78003 87141
rect 79200 87138 80000 87168
rect 77937 87136 80000 87138
rect 77937 87080 77942 87136
rect 77998 87080 80000 87136
rect 77937 87078 80000 87080
rect 77937 87075 78003 87078
rect 19568 87072 19888 87073
rect 19568 87008 19576 87072
rect 19640 87008 19656 87072
rect 19720 87008 19736 87072
rect 19800 87008 19816 87072
rect 19880 87008 19888 87072
rect 19568 87007 19888 87008
rect 50288 87072 50608 87073
rect 50288 87008 50296 87072
rect 50360 87008 50376 87072
rect 50440 87008 50456 87072
rect 50520 87008 50536 87072
rect 50600 87008 50608 87072
rect 79200 87048 80000 87078
rect 50288 87007 50608 87008
rect 4208 86528 4528 86529
rect 4208 86464 4216 86528
rect 4280 86464 4296 86528
rect 4360 86464 4376 86528
rect 4440 86464 4456 86528
rect 4520 86464 4528 86528
rect 4208 86463 4528 86464
rect 34928 86528 35248 86529
rect 34928 86464 34936 86528
rect 35000 86464 35016 86528
rect 35080 86464 35096 86528
rect 35160 86464 35176 86528
rect 35240 86464 35248 86528
rect 34928 86463 35248 86464
rect 65648 86528 65968 86529
rect 65648 86464 65656 86528
rect 65720 86464 65736 86528
rect 65800 86464 65816 86528
rect 65880 86464 65896 86528
rect 65960 86464 65968 86528
rect 65648 86463 65968 86464
rect 19568 85984 19888 85985
rect 19568 85920 19576 85984
rect 19640 85920 19656 85984
rect 19720 85920 19736 85984
rect 19800 85920 19816 85984
rect 19880 85920 19888 85984
rect 19568 85919 19888 85920
rect 50288 85984 50608 85985
rect 50288 85920 50296 85984
rect 50360 85920 50376 85984
rect 50440 85920 50456 85984
rect 50520 85920 50536 85984
rect 50600 85920 50608 85984
rect 50288 85919 50608 85920
rect 0 85778 800 85808
rect 1577 85778 1643 85781
rect 0 85776 1643 85778
rect 0 85720 1582 85776
rect 1638 85720 1643 85776
rect 0 85718 1643 85720
rect 0 85688 800 85718
rect 1577 85715 1643 85718
rect 4208 85440 4528 85441
rect 4208 85376 4216 85440
rect 4280 85376 4296 85440
rect 4360 85376 4376 85440
rect 4440 85376 4456 85440
rect 4520 85376 4528 85440
rect 4208 85375 4528 85376
rect 34928 85440 35248 85441
rect 34928 85376 34936 85440
rect 35000 85376 35016 85440
rect 35080 85376 35096 85440
rect 35160 85376 35176 85440
rect 35240 85376 35248 85440
rect 34928 85375 35248 85376
rect 65648 85440 65968 85441
rect 65648 85376 65656 85440
rect 65720 85376 65736 85440
rect 65800 85376 65816 85440
rect 65880 85376 65896 85440
rect 65960 85376 65968 85440
rect 65648 85375 65968 85376
rect 19568 84896 19888 84897
rect 19568 84832 19576 84896
rect 19640 84832 19656 84896
rect 19720 84832 19736 84896
rect 19800 84832 19816 84896
rect 19880 84832 19888 84896
rect 19568 84831 19888 84832
rect 50288 84896 50608 84897
rect 50288 84832 50296 84896
rect 50360 84832 50376 84896
rect 50440 84832 50456 84896
rect 50520 84832 50536 84896
rect 50600 84832 50608 84896
rect 50288 84831 50608 84832
rect 4208 84352 4528 84353
rect 4208 84288 4216 84352
rect 4280 84288 4296 84352
rect 4360 84288 4376 84352
rect 4440 84288 4456 84352
rect 4520 84288 4528 84352
rect 4208 84287 4528 84288
rect 34928 84352 35248 84353
rect 34928 84288 34936 84352
rect 35000 84288 35016 84352
rect 35080 84288 35096 84352
rect 35160 84288 35176 84352
rect 35240 84288 35248 84352
rect 34928 84287 35248 84288
rect 65648 84352 65968 84353
rect 65648 84288 65656 84352
rect 65720 84288 65736 84352
rect 65800 84288 65816 84352
rect 65880 84288 65896 84352
rect 65960 84288 65968 84352
rect 65648 84287 65968 84288
rect 19568 83808 19888 83809
rect 19568 83744 19576 83808
rect 19640 83744 19656 83808
rect 19720 83744 19736 83808
rect 19800 83744 19816 83808
rect 19880 83744 19888 83808
rect 19568 83743 19888 83744
rect 50288 83808 50608 83809
rect 50288 83744 50296 83808
rect 50360 83744 50376 83808
rect 50440 83744 50456 83808
rect 50520 83744 50536 83808
rect 50600 83744 50608 83808
rect 50288 83743 50608 83744
rect 4208 83264 4528 83265
rect 4208 83200 4216 83264
rect 4280 83200 4296 83264
rect 4360 83200 4376 83264
rect 4440 83200 4456 83264
rect 4520 83200 4528 83264
rect 4208 83199 4528 83200
rect 34928 83264 35248 83265
rect 34928 83200 34936 83264
rect 35000 83200 35016 83264
rect 35080 83200 35096 83264
rect 35160 83200 35176 83264
rect 35240 83200 35248 83264
rect 34928 83199 35248 83200
rect 65648 83264 65968 83265
rect 65648 83200 65656 83264
rect 65720 83200 65736 83264
rect 65800 83200 65816 83264
rect 65880 83200 65896 83264
rect 65960 83200 65968 83264
rect 65648 83199 65968 83200
rect 77845 83058 77911 83061
rect 79200 83058 80000 83088
rect 77845 83056 80000 83058
rect 77845 83000 77850 83056
rect 77906 83000 80000 83056
rect 77845 82998 80000 83000
rect 77845 82995 77911 82998
rect 79200 82968 80000 82998
rect 19568 82720 19888 82721
rect 19568 82656 19576 82720
rect 19640 82656 19656 82720
rect 19720 82656 19736 82720
rect 19800 82656 19816 82720
rect 19880 82656 19888 82720
rect 19568 82655 19888 82656
rect 50288 82720 50608 82721
rect 50288 82656 50296 82720
rect 50360 82656 50376 82720
rect 50440 82656 50456 82720
rect 50520 82656 50536 82720
rect 50600 82656 50608 82720
rect 50288 82655 50608 82656
rect 4208 82176 4528 82177
rect 4208 82112 4216 82176
rect 4280 82112 4296 82176
rect 4360 82112 4376 82176
rect 4440 82112 4456 82176
rect 4520 82112 4528 82176
rect 4208 82111 4528 82112
rect 34928 82176 35248 82177
rect 34928 82112 34936 82176
rect 35000 82112 35016 82176
rect 35080 82112 35096 82176
rect 35160 82112 35176 82176
rect 35240 82112 35248 82176
rect 34928 82111 35248 82112
rect 65648 82176 65968 82177
rect 65648 82112 65656 82176
rect 65720 82112 65736 82176
rect 65800 82112 65816 82176
rect 65880 82112 65896 82176
rect 65960 82112 65968 82176
rect 65648 82111 65968 82112
rect 0 81698 800 81728
rect 1393 81698 1459 81701
rect 0 81696 1459 81698
rect 0 81640 1398 81696
rect 1454 81640 1459 81696
rect 0 81638 1459 81640
rect 0 81608 800 81638
rect 1393 81635 1459 81638
rect 19568 81632 19888 81633
rect 19568 81568 19576 81632
rect 19640 81568 19656 81632
rect 19720 81568 19736 81632
rect 19800 81568 19816 81632
rect 19880 81568 19888 81632
rect 19568 81567 19888 81568
rect 50288 81632 50608 81633
rect 50288 81568 50296 81632
rect 50360 81568 50376 81632
rect 50440 81568 50456 81632
rect 50520 81568 50536 81632
rect 50600 81568 50608 81632
rect 50288 81567 50608 81568
rect 4208 81088 4528 81089
rect 4208 81024 4216 81088
rect 4280 81024 4296 81088
rect 4360 81024 4376 81088
rect 4440 81024 4456 81088
rect 4520 81024 4528 81088
rect 4208 81023 4528 81024
rect 34928 81088 35248 81089
rect 34928 81024 34936 81088
rect 35000 81024 35016 81088
rect 35080 81024 35096 81088
rect 35160 81024 35176 81088
rect 35240 81024 35248 81088
rect 34928 81023 35248 81024
rect 65648 81088 65968 81089
rect 65648 81024 65656 81088
rect 65720 81024 65736 81088
rect 65800 81024 65816 81088
rect 65880 81024 65896 81088
rect 65960 81024 65968 81088
rect 65648 81023 65968 81024
rect 19568 80544 19888 80545
rect 19568 80480 19576 80544
rect 19640 80480 19656 80544
rect 19720 80480 19736 80544
rect 19800 80480 19816 80544
rect 19880 80480 19888 80544
rect 19568 80479 19888 80480
rect 50288 80544 50608 80545
rect 50288 80480 50296 80544
rect 50360 80480 50376 80544
rect 50440 80480 50456 80544
rect 50520 80480 50536 80544
rect 50600 80480 50608 80544
rect 50288 80479 50608 80480
rect 4208 80000 4528 80001
rect 4208 79936 4216 80000
rect 4280 79936 4296 80000
rect 4360 79936 4376 80000
rect 4440 79936 4456 80000
rect 4520 79936 4528 80000
rect 4208 79935 4528 79936
rect 34928 80000 35248 80001
rect 34928 79936 34936 80000
rect 35000 79936 35016 80000
rect 35080 79936 35096 80000
rect 35160 79936 35176 80000
rect 35240 79936 35248 80000
rect 34928 79935 35248 79936
rect 65648 80000 65968 80001
rect 65648 79936 65656 80000
rect 65720 79936 65736 80000
rect 65800 79936 65816 80000
rect 65880 79936 65896 80000
rect 65960 79936 65968 80000
rect 65648 79935 65968 79936
rect 19568 79456 19888 79457
rect 19568 79392 19576 79456
rect 19640 79392 19656 79456
rect 19720 79392 19736 79456
rect 19800 79392 19816 79456
rect 19880 79392 19888 79456
rect 19568 79391 19888 79392
rect 50288 79456 50608 79457
rect 50288 79392 50296 79456
rect 50360 79392 50376 79456
rect 50440 79392 50456 79456
rect 50520 79392 50536 79456
rect 50600 79392 50608 79456
rect 50288 79391 50608 79392
rect 77569 78978 77635 78981
rect 79200 78978 80000 79008
rect 77569 78976 80000 78978
rect 77569 78920 77574 78976
rect 77630 78920 80000 78976
rect 77569 78918 80000 78920
rect 77569 78915 77635 78918
rect 4208 78912 4528 78913
rect 4208 78848 4216 78912
rect 4280 78848 4296 78912
rect 4360 78848 4376 78912
rect 4440 78848 4456 78912
rect 4520 78848 4528 78912
rect 4208 78847 4528 78848
rect 34928 78912 35248 78913
rect 34928 78848 34936 78912
rect 35000 78848 35016 78912
rect 35080 78848 35096 78912
rect 35160 78848 35176 78912
rect 35240 78848 35248 78912
rect 34928 78847 35248 78848
rect 65648 78912 65968 78913
rect 65648 78848 65656 78912
rect 65720 78848 65736 78912
rect 65800 78848 65816 78912
rect 65880 78848 65896 78912
rect 65960 78848 65968 78912
rect 79200 78888 80000 78918
rect 65648 78847 65968 78848
rect 19568 78368 19888 78369
rect 0 78298 800 78328
rect 19568 78304 19576 78368
rect 19640 78304 19656 78368
rect 19720 78304 19736 78368
rect 19800 78304 19816 78368
rect 19880 78304 19888 78368
rect 19568 78303 19888 78304
rect 50288 78368 50608 78369
rect 50288 78304 50296 78368
rect 50360 78304 50376 78368
rect 50440 78304 50456 78368
rect 50520 78304 50536 78368
rect 50600 78304 50608 78368
rect 50288 78303 50608 78304
rect 1577 78298 1643 78301
rect 0 78296 1643 78298
rect 0 78240 1582 78296
rect 1638 78240 1643 78296
rect 0 78238 1643 78240
rect 0 78208 800 78238
rect 1577 78235 1643 78238
rect 4208 77824 4528 77825
rect 4208 77760 4216 77824
rect 4280 77760 4296 77824
rect 4360 77760 4376 77824
rect 4440 77760 4456 77824
rect 4520 77760 4528 77824
rect 4208 77759 4528 77760
rect 34928 77824 35248 77825
rect 34928 77760 34936 77824
rect 35000 77760 35016 77824
rect 35080 77760 35096 77824
rect 35160 77760 35176 77824
rect 35240 77760 35248 77824
rect 34928 77759 35248 77760
rect 65648 77824 65968 77825
rect 65648 77760 65656 77824
rect 65720 77760 65736 77824
rect 65800 77760 65816 77824
rect 65880 77760 65896 77824
rect 65960 77760 65968 77824
rect 65648 77759 65968 77760
rect 19568 77280 19888 77281
rect 19568 77216 19576 77280
rect 19640 77216 19656 77280
rect 19720 77216 19736 77280
rect 19800 77216 19816 77280
rect 19880 77216 19888 77280
rect 19568 77215 19888 77216
rect 50288 77280 50608 77281
rect 50288 77216 50296 77280
rect 50360 77216 50376 77280
rect 50440 77216 50456 77280
rect 50520 77216 50536 77280
rect 50600 77216 50608 77280
rect 50288 77215 50608 77216
rect 4208 76736 4528 76737
rect 4208 76672 4216 76736
rect 4280 76672 4296 76736
rect 4360 76672 4376 76736
rect 4440 76672 4456 76736
rect 4520 76672 4528 76736
rect 4208 76671 4528 76672
rect 34928 76736 35248 76737
rect 34928 76672 34936 76736
rect 35000 76672 35016 76736
rect 35080 76672 35096 76736
rect 35160 76672 35176 76736
rect 35240 76672 35248 76736
rect 34928 76671 35248 76672
rect 65648 76736 65968 76737
rect 65648 76672 65656 76736
rect 65720 76672 65736 76736
rect 65800 76672 65816 76736
rect 65880 76672 65896 76736
rect 65960 76672 65968 76736
rect 65648 76671 65968 76672
rect 19568 76192 19888 76193
rect 19568 76128 19576 76192
rect 19640 76128 19656 76192
rect 19720 76128 19736 76192
rect 19800 76128 19816 76192
rect 19880 76128 19888 76192
rect 19568 76127 19888 76128
rect 50288 76192 50608 76193
rect 50288 76128 50296 76192
rect 50360 76128 50376 76192
rect 50440 76128 50456 76192
rect 50520 76128 50536 76192
rect 50600 76128 50608 76192
rect 50288 76127 50608 76128
rect 4208 75648 4528 75649
rect 4208 75584 4216 75648
rect 4280 75584 4296 75648
rect 4360 75584 4376 75648
rect 4440 75584 4456 75648
rect 4520 75584 4528 75648
rect 4208 75583 4528 75584
rect 34928 75648 35248 75649
rect 34928 75584 34936 75648
rect 35000 75584 35016 75648
rect 35080 75584 35096 75648
rect 35160 75584 35176 75648
rect 35240 75584 35248 75648
rect 34928 75583 35248 75584
rect 65648 75648 65968 75649
rect 65648 75584 65656 75648
rect 65720 75584 65736 75648
rect 65800 75584 65816 75648
rect 65880 75584 65896 75648
rect 65960 75584 65968 75648
rect 65648 75583 65968 75584
rect 19568 75104 19888 75105
rect 19568 75040 19576 75104
rect 19640 75040 19656 75104
rect 19720 75040 19736 75104
rect 19800 75040 19816 75104
rect 19880 75040 19888 75104
rect 19568 75039 19888 75040
rect 50288 75104 50608 75105
rect 50288 75040 50296 75104
rect 50360 75040 50376 75104
rect 50440 75040 50456 75104
rect 50520 75040 50536 75104
rect 50600 75040 50608 75104
rect 50288 75039 50608 75040
rect 78029 74898 78095 74901
rect 79200 74898 80000 74928
rect 78029 74896 80000 74898
rect 78029 74840 78034 74896
rect 78090 74840 80000 74896
rect 78029 74838 80000 74840
rect 78029 74835 78095 74838
rect 79200 74808 80000 74838
rect 4208 74560 4528 74561
rect 4208 74496 4216 74560
rect 4280 74496 4296 74560
rect 4360 74496 4376 74560
rect 4440 74496 4456 74560
rect 4520 74496 4528 74560
rect 4208 74495 4528 74496
rect 34928 74560 35248 74561
rect 34928 74496 34936 74560
rect 35000 74496 35016 74560
rect 35080 74496 35096 74560
rect 35160 74496 35176 74560
rect 35240 74496 35248 74560
rect 34928 74495 35248 74496
rect 65648 74560 65968 74561
rect 65648 74496 65656 74560
rect 65720 74496 65736 74560
rect 65800 74496 65816 74560
rect 65880 74496 65896 74560
rect 65960 74496 65968 74560
rect 65648 74495 65968 74496
rect 0 74218 800 74248
rect 1577 74218 1643 74221
rect 0 74216 1643 74218
rect 0 74160 1582 74216
rect 1638 74160 1643 74216
rect 0 74158 1643 74160
rect 0 74128 800 74158
rect 1577 74155 1643 74158
rect 19568 74016 19888 74017
rect 19568 73952 19576 74016
rect 19640 73952 19656 74016
rect 19720 73952 19736 74016
rect 19800 73952 19816 74016
rect 19880 73952 19888 74016
rect 19568 73951 19888 73952
rect 50288 74016 50608 74017
rect 50288 73952 50296 74016
rect 50360 73952 50376 74016
rect 50440 73952 50456 74016
rect 50520 73952 50536 74016
rect 50600 73952 50608 74016
rect 50288 73951 50608 73952
rect 4208 73472 4528 73473
rect 4208 73408 4216 73472
rect 4280 73408 4296 73472
rect 4360 73408 4376 73472
rect 4440 73408 4456 73472
rect 4520 73408 4528 73472
rect 4208 73407 4528 73408
rect 34928 73472 35248 73473
rect 34928 73408 34936 73472
rect 35000 73408 35016 73472
rect 35080 73408 35096 73472
rect 35160 73408 35176 73472
rect 35240 73408 35248 73472
rect 34928 73407 35248 73408
rect 65648 73472 65968 73473
rect 65648 73408 65656 73472
rect 65720 73408 65736 73472
rect 65800 73408 65816 73472
rect 65880 73408 65896 73472
rect 65960 73408 65968 73472
rect 65648 73407 65968 73408
rect 19568 72928 19888 72929
rect 19568 72864 19576 72928
rect 19640 72864 19656 72928
rect 19720 72864 19736 72928
rect 19800 72864 19816 72928
rect 19880 72864 19888 72928
rect 19568 72863 19888 72864
rect 50288 72928 50608 72929
rect 50288 72864 50296 72928
rect 50360 72864 50376 72928
rect 50440 72864 50456 72928
rect 50520 72864 50536 72928
rect 50600 72864 50608 72928
rect 50288 72863 50608 72864
rect 4208 72384 4528 72385
rect 4208 72320 4216 72384
rect 4280 72320 4296 72384
rect 4360 72320 4376 72384
rect 4440 72320 4456 72384
rect 4520 72320 4528 72384
rect 4208 72319 4528 72320
rect 34928 72384 35248 72385
rect 34928 72320 34936 72384
rect 35000 72320 35016 72384
rect 35080 72320 35096 72384
rect 35160 72320 35176 72384
rect 35240 72320 35248 72384
rect 34928 72319 35248 72320
rect 65648 72384 65968 72385
rect 65648 72320 65656 72384
rect 65720 72320 65736 72384
rect 65800 72320 65816 72384
rect 65880 72320 65896 72384
rect 65960 72320 65968 72384
rect 65648 72319 65968 72320
rect 19568 71840 19888 71841
rect 19568 71776 19576 71840
rect 19640 71776 19656 71840
rect 19720 71776 19736 71840
rect 19800 71776 19816 71840
rect 19880 71776 19888 71840
rect 19568 71775 19888 71776
rect 50288 71840 50608 71841
rect 50288 71776 50296 71840
rect 50360 71776 50376 71840
rect 50440 71776 50456 71840
rect 50520 71776 50536 71840
rect 50600 71776 50608 71840
rect 50288 71775 50608 71776
rect 77845 71498 77911 71501
rect 79200 71498 80000 71528
rect 77845 71496 80000 71498
rect 77845 71440 77850 71496
rect 77906 71440 80000 71496
rect 77845 71438 80000 71440
rect 77845 71435 77911 71438
rect 79200 71408 80000 71438
rect 4208 71296 4528 71297
rect 4208 71232 4216 71296
rect 4280 71232 4296 71296
rect 4360 71232 4376 71296
rect 4440 71232 4456 71296
rect 4520 71232 4528 71296
rect 4208 71231 4528 71232
rect 34928 71296 35248 71297
rect 34928 71232 34936 71296
rect 35000 71232 35016 71296
rect 35080 71232 35096 71296
rect 35160 71232 35176 71296
rect 35240 71232 35248 71296
rect 34928 71231 35248 71232
rect 65648 71296 65968 71297
rect 65648 71232 65656 71296
rect 65720 71232 65736 71296
rect 65800 71232 65816 71296
rect 65880 71232 65896 71296
rect 65960 71232 65968 71296
rect 65648 71231 65968 71232
rect 19568 70752 19888 70753
rect 19568 70688 19576 70752
rect 19640 70688 19656 70752
rect 19720 70688 19736 70752
rect 19800 70688 19816 70752
rect 19880 70688 19888 70752
rect 19568 70687 19888 70688
rect 50288 70752 50608 70753
rect 50288 70688 50296 70752
rect 50360 70688 50376 70752
rect 50440 70688 50456 70752
rect 50520 70688 50536 70752
rect 50600 70688 50608 70752
rect 50288 70687 50608 70688
rect 4208 70208 4528 70209
rect 0 70138 800 70168
rect 4208 70144 4216 70208
rect 4280 70144 4296 70208
rect 4360 70144 4376 70208
rect 4440 70144 4456 70208
rect 4520 70144 4528 70208
rect 4208 70143 4528 70144
rect 34928 70208 35248 70209
rect 34928 70144 34936 70208
rect 35000 70144 35016 70208
rect 35080 70144 35096 70208
rect 35160 70144 35176 70208
rect 35240 70144 35248 70208
rect 34928 70143 35248 70144
rect 65648 70208 65968 70209
rect 65648 70144 65656 70208
rect 65720 70144 65736 70208
rect 65800 70144 65816 70208
rect 65880 70144 65896 70208
rect 65960 70144 65968 70208
rect 65648 70143 65968 70144
rect 1577 70138 1643 70141
rect 0 70136 1643 70138
rect 0 70080 1582 70136
rect 1638 70080 1643 70136
rect 0 70078 1643 70080
rect 0 70048 800 70078
rect 1577 70075 1643 70078
rect 19568 69664 19888 69665
rect 19568 69600 19576 69664
rect 19640 69600 19656 69664
rect 19720 69600 19736 69664
rect 19800 69600 19816 69664
rect 19880 69600 19888 69664
rect 19568 69599 19888 69600
rect 50288 69664 50608 69665
rect 50288 69600 50296 69664
rect 50360 69600 50376 69664
rect 50440 69600 50456 69664
rect 50520 69600 50536 69664
rect 50600 69600 50608 69664
rect 50288 69599 50608 69600
rect 4208 69120 4528 69121
rect 4208 69056 4216 69120
rect 4280 69056 4296 69120
rect 4360 69056 4376 69120
rect 4440 69056 4456 69120
rect 4520 69056 4528 69120
rect 4208 69055 4528 69056
rect 34928 69120 35248 69121
rect 34928 69056 34936 69120
rect 35000 69056 35016 69120
rect 35080 69056 35096 69120
rect 35160 69056 35176 69120
rect 35240 69056 35248 69120
rect 34928 69055 35248 69056
rect 65648 69120 65968 69121
rect 65648 69056 65656 69120
rect 65720 69056 65736 69120
rect 65800 69056 65816 69120
rect 65880 69056 65896 69120
rect 65960 69056 65968 69120
rect 65648 69055 65968 69056
rect 19568 68576 19888 68577
rect 19568 68512 19576 68576
rect 19640 68512 19656 68576
rect 19720 68512 19736 68576
rect 19800 68512 19816 68576
rect 19880 68512 19888 68576
rect 19568 68511 19888 68512
rect 50288 68576 50608 68577
rect 50288 68512 50296 68576
rect 50360 68512 50376 68576
rect 50440 68512 50456 68576
rect 50520 68512 50536 68576
rect 50600 68512 50608 68576
rect 50288 68511 50608 68512
rect 4208 68032 4528 68033
rect 4208 67968 4216 68032
rect 4280 67968 4296 68032
rect 4360 67968 4376 68032
rect 4440 67968 4456 68032
rect 4520 67968 4528 68032
rect 4208 67967 4528 67968
rect 34928 68032 35248 68033
rect 34928 67968 34936 68032
rect 35000 67968 35016 68032
rect 35080 67968 35096 68032
rect 35160 67968 35176 68032
rect 35240 67968 35248 68032
rect 34928 67967 35248 67968
rect 65648 68032 65968 68033
rect 65648 67968 65656 68032
rect 65720 67968 65736 68032
rect 65800 67968 65816 68032
rect 65880 67968 65896 68032
rect 65960 67968 65968 68032
rect 65648 67967 65968 67968
rect 19568 67488 19888 67489
rect 19568 67424 19576 67488
rect 19640 67424 19656 67488
rect 19720 67424 19736 67488
rect 19800 67424 19816 67488
rect 19880 67424 19888 67488
rect 19568 67423 19888 67424
rect 50288 67488 50608 67489
rect 50288 67424 50296 67488
rect 50360 67424 50376 67488
rect 50440 67424 50456 67488
rect 50520 67424 50536 67488
rect 50600 67424 50608 67488
rect 50288 67423 50608 67424
rect 77937 67418 78003 67421
rect 79200 67418 80000 67448
rect 77937 67416 80000 67418
rect 77937 67360 77942 67416
rect 77998 67360 80000 67416
rect 77937 67358 80000 67360
rect 77937 67355 78003 67358
rect 79200 67328 80000 67358
rect 4208 66944 4528 66945
rect 4208 66880 4216 66944
rect 4280 66880 4296 66944
rect 4360 66880 4376 66944
rect 4440 66880 4456 66944
rect 4520 66880 4528 66944
rect 4208 66879 4528 66880
rect 34928 66944 35248 66945
rect 34928 66880 34936 66944
rect 35000 66880 35016 66944
rect 35080 66880 35096 66944
rect 35160 66880 35176 66944
rect 35240 66880 35248 66944
rect 34928 66879 35248 66880
rect 65648 66944 65968 66945
rect 65648 66880 65656 66944
rect 65720 66880 65736 66944
rect 65800 66880 65816 66944
rect 65880 66880 65896 66944
rect 65960 66880 65968 66944
rect 65648 66879 65968 66880
rect 19568 66400 19888 66401
rect 19568 66336 19576 66400
rect 19640 66336 19656 66400
rect 19720 66336 19736 66400
rect 19800 66336 19816 66400
rect 19880 66336 19888 66400
rect 19568 66335 19888 66336
rect 50288 66400 50608 66401
rect 50288 66336 50296 66400
rect 50360 66336 50376 66400
rect 50440 66336 50456 66400
rect 50520 66336 50536 66400
rect 50600 66336 50608 66400
rect 50288 66335 50608 66336
rect 0 66058 800 66088
rect 1577 66058 1643 66061
rect 0 66056 1643 66058
rect 0 66000 1582 66056
rect 1638 66000 1643 66056
rect 0 65998 1643 66000
rect 0 65968 800 65998
rect 1577 65995 1643 65998
rect 4208 65856 4528 65857
rect 4208 65792 4216 65856
rect 4280 65792 4296 65856
rect 4360 65792 4376 65856
rect 4440 65792 4456 65856
rect 4520 65792 4528 65856
rect 4208 65791 4528 65792
rect 34928 65856 35248 65857
rect 34928 65792 34936 65856
rect 35000 65792 35016 65856
rect 35080 65792 35096 65856
rect 35160 65792 35176 65856
rect 35240 65792 35248 65856
rect 34928 65791 35248 65792
rect 65648 65856 65968 65857
rect 65648 65792 65656 65856
rect 65720 65792 65736 65856
rect 65800 65792 65816 65856
rect 65880 65792 65896 65856
rect 65960 65792 65968 65856
rect 65648 65791 65968 65792
rect 19568 65312 19888 65313
rect 19568 65248 19576 65312
rect 19640 65248 19656 65312
rect 19720 65248 19736 65312
rect 19800 65248 19816 65312
rect 19880 65248 19888 65312
rect 19568 65247 19888 65248
rect 50288 65312 50608 65313
rect 50288 65248 50296 65312
rect 50360 65248 50376 65312
rect 50440 65248 50456 65312
rect 50520 65248 50536 65312
rect 50600 65248 50608 65312
rect 50288 65247 50608 65248
rect 4208 64768 4528 64769
rect 4208 64704 4216 64768
rect 4280 64704 4296 64768
rect 4360 64704 4376 64768
rect 4440 64704 4456 64768
rect 4520 64704 4528 64768
rect 4208 64703 4528 64704
rect 34928 64768 35248 64769
rect 34928 64704 34936 64768
rect 35000 64704 35016 64768
rect 35080 64704 35096 64768
rect 35160 64704 35176 64768
rect 35240 64704 35248 64768
rect 34928 64703 35248 64704
rect 65648 64768 65968 64769
rect 65648 64704 65656 64768
rect 65720 64704 65736 64768
rect 65800 64704 65816 64768
rect 65880 64704 65896 64768
rect 65960 64704 65968 64768
rect 65648 64703 65968 64704
rect 19568 64224 19888 64225
rect 19568 64160 19576 64224
rect 19640 64160 19656 64224
rect 19720 64160 19736 64224
rect 19800 64160 19816 64224
rect 19880 64160 19888 64224
rect 19568 64159 19888 64160
rect 50288 64224 50608 64225
rect 50288 64160 50296 64224
rect 50360 64160 50376 64224
rect 50440 64160 50456 64224
rect 50520 64160 50536 64224
rect 50600 64160 50608 64224
rect 50288 64159 50608 64160
rect 4208 63680 4528 63681
rect 4208 63616 4216 63680
rect 4280 63616 4296 63680
rect 4360 63616 4376 63680
rect 4440 63616 4456 63680
rect 4520 63616 4528 63680
rect 4208 63615 4528 63616
rect 34928 63680 35248 63681
rect 34928 63616 34936 63680
rect 35000 63616 35016 63680
rect 35080 63616 35096 63680
rect 35160 63616 35176 63680
rect 35240 63616 35248 63680
rect 34928 63615 35248 63616
rect 65648 63680 65968 63681
rect 65648 63616 65656 63680
rect 65720 63616 65736 63680
rect 65800 63616 65816 63680
rect 65880 63616 65896 63680
rect 65960 63616 65968 63680
rect 65648 63615 65968 63616
rect 78029 63338 78095 63341
rect 79200 63338 80000 63368
rect 78029 63336 80000 63338
rect 78029 63280 78034 63336
rect 78090 63280 80000 63336
rect 78029 63278 80000 63280
rect 78029 63275 78095 63278
rect 79200 63248 80000 63278
rect 19568 63136 19888 63137
rect 19568 63072 19576 63136
rect 19640 63072 19656 63136
rect 19720 63072 19736 63136
rect 19800 63072 19816 63136
rect 19880 63072 19888 63136
rect 19568 63071 19888 63072
rect 50288 63136 50608 63137
rect 50288 63072 50296 63136
rect 50360 63072 50376 63136
rect 50440 63072 50456 63136
rect 50520 63072 50536 63136
rect 50600 63072 50608 63136
rect 50288 63071 50608 63072
rect 0 62658 800 62688
rect 1577 62658 1643 62661
rect 0 62656 1643 62658
rect 0 62600 1582 62656
rect 1638 62600 1643 62656
rect 0 62598 1643 62600
rect 0 62568 800 62598
rect 1577 62595 1643 62598
rect 4208 62592 4528 62593
rect 4208 62528 4216 62592
rect 4280 62528 4296 62592
rect 4360 62528 4376 62592
rect 4440 62528 4456 62592
rect 4520 62528 4528 62592
rect 4208 62527 4528 62528
rect 34928 62592 35248 62593
rect 34928 62528 34936 62592
rect 35000 62528 35016 62592
rect 35080 62528 35096 62592
rect 35160 62528 35176 62592
rect 35240 62528 35248 62592
rect 34928 62527 35248 62528
rect 65648 62592 65968 62593
rect 65648 62528 65656 62592
rect 65720 62528 65736 62592
rect 65800 62528 65816 62592
rect 65880 62528 65896 62592
rect 65960 62528 65968 62592
rect 65648 62527 65968 62528
rect 19568 62048 19888 62049
rect 19568 61984 19576 62048
rect 19640 61984 19656 62048
rect 19720 61984 19736 62048
rect 19800 61984 19816 62048
rect 19880 61984 19888 62048
rect 19568 61983 19888 61984
rect 50288 62048 50608 62049
rect 50288 61984 50296 62048
rect 50360 61984 50376 62048
rect 50440 61984 50456 62048
rect 50520 61984 50536 62048
rect 50600 61984 50608 62048
rect 50288 61983 50608 61984
rect 4208 61504 4528 61505
rect 4208 61440 4216 61504
rect 4280 61440 4296 61504
rect 4360 61440 4376 61504
rect 4440 61440 4456 61504
rect 4520 61440 4528 61504
rect 4208 61439 4528 61440
rect 34928 61504 35248 61505
rect 34928 61440 34936 61504
rect 35000 61440 35016 61504
rect 35080 61440 35096 61504
rect 35160 61440 35176 61504
rect 35240 61440 35248 61504
rect 34928 61439 35248 61440
rect 65648 61504 65968 61505
rect 65648 61440 65656 61504
rect 65720 61440 65736 61504
rect 65800 61440 65816 61504
rect 65880 61440 65896 61504
rect 65960 61440 65968 61504
rect 65648 61439 65968 61440
rect 19568 60960 19888 60961
rect 19568 60896 19576 60960
rect 19640 60896 19656 60960
rect 19720 60896 19736 60960
rect 19800 60896 19816 60960
rect 19880 60896 19888 60960
rect 19568 60895 19888 60896
rect 50288 60960 50608 60961
rect 50288 60896 50296 60960
rect 50360 60896 50376 60960
rect 50440 60896 50456 60960
rect 50520 60896 50536 60960
rect 50600 60896 50608 60960
rect 50288 60895 50608 60896
rect 4208 60416 4528 60417
rect 4208 60352 4216 60416
rect 4280 60352 4296 60416
rect 4360 60352 4376 60416
rect 4440 60352 4456 60416
rect 4520 60352 4528 60416
rect 4208 60351 4528 60352
rect 34928 60416 35248 60417
rect 34928 60352 34936 60416
rect 35000 60352 35016 60416
rect 35080 60352 35096 60416
rect 35160 60352 35176 60416
rect 35240 60352 35248 60416
rect 34928 60351 35248 60352
rect 65648 60416 65968 60417
rect 65648 60352 65656 60416
rect 65720 60352 65736 60416
rect 65800 60352 65816 60416
rect 65880 60352 65896 60416
rect 65960 60352 65968 60416
rect 65648 60351 65968 60352
rect 19568 59872 19888 59873
rect 19568 59808 19576 59872
rect 19640 59808 19656 59872
rect 19720 59808 19736 59872
rect 19800 59808 19816 59872
rect 19880 59808 19888 59872
rect 19568 59807 19888 59808
rect 50288 59872 50608 59873
rect 50288 59808 50296 59872
rect 50360 59808 50376 59872
rect 50440 59808 50456 59872
rect 50520 59808 50536 59872
rect 50600 59808 50608 59872
rect 50288 59807 50608 59808
rect 4208 59328 4528 59329
rect 4208 59264 4216 59328
rect 4280 59264 4296 59328
rect 4360 59264 4376 59328
rect 4440 59264 4456 59328
rect 4520 59264 4528 59328
rect 4208 59263 4528 59264
rect 34928 59328 35248 59329
rect 34928 59264 34936 59328
rect 35000 59264 35016 59328
rect 35080 59264 35096 59328
rect 35160 59264 35176 59328
rect 35240 59264 35248 59328
rect 34928 59263 35248 59264
rect 65648 59328 65968 59329
rect 65648 59264 65656 59328
rect 65720 59264 65736 59328
rect 65800 59264 65816 59328
rect 65880 59264 65896 59328
rect 65960 59264 65968 59328
rect 65648 59263 65968 59264
rect 77937 59258 78003 59261
rect 79200 59258 80000 59288
rect 77937 59256 80000 59258
rect 77937 59200 77942 59256
rect 77998 59200 80000 59256
rect 77937 59198 80000 59200
rect 77937 59195 78003 59198
rect 79200 59168 80000 59198
rect 19568 58784 19888 58785
rect 19568 58720 19576 58784
rect 19640 58720 19656 58784
rect 19720 58720 19736 58784
rect 19800 58720 19816 58784
rect 19880 58720 19888 58784
rect 19568 58719 19888 58720
rect 50288 58784 50608 58785
rect 50288 58720 50296 58784
rect 50360 58720 50376 58784
rect 50440 58720 50456 58784
rect 50520 58720 50536 58784
rect 50600 58720 50608 58784
rect 50288 58719 50608 58720
rect 0 58578 800 58608
rect 1577 58578 1643 58581
rect 0 58576 1643 58578
rect 0 58520 1582 58576
rect 1638 58520 1643 58576
rect 0 58518 1643 58520
rect 0 58488 800 58518
rect 1577 58515 1643 58518
rect 4208 58240 4528 58241
rect 4208 58176 4216 58240
rect 4280 58176 4296 58240
rect 4360 58176 4376 58240
rect 4440 58176 4456 58240
rect 4520 58176 4528 58240
rect 4208 58175 4528 58176
rect 34928 58240 35248 58241
rect 34928 58176 34936 58240
rect 35000 58176 35016 58240
rect 35080 58176 35096 58240
rect 35160 58176 35176 58240
rect 35240 58176 35248 58240
rect 34928 58175 35248 58176
rect 65648 58240 65968 58241
rect 65648 58176 65656 58240
rect 65720 58176 65736 58240
rect 65800 58176 65816 58240
rect 65880 58176 65896 58240
rect 65960 58176 65968 58240
rect 65648 58175 65968 58176
rect 19568 57696 19888 57697
rect 19568 57632 19576 57696
rect 19640 57632 19656 57696
rect 19720 57632 19736 57696
rect 19800 57632 19816 57696
rect 19880 57632 19888 57696
rect 19568 57631 19888 57632
rect 50288 57696 50608 57697
rect 50288 57632 50296 57696
rect 50360 57632 50376 57696
rect 50440 57632 50456 57696
rect 50520 57632 50536 57696
rect 50600 57632 50608 57696
rect 50288 57631 50608 57632
rect 4208 57152 4528 57153
rect 4208 57088 4216 57152
rect 4280 57088 4296 57152
rect 4360 57088 4376 57152
rect 4440 57088 4456 57152
rect 4520 57088 4528 57152
rect 4208 57087 4528 57088
rect 34928 57152 35248 57153
rect 34928 57088 34936 57152
rect 35000 57088 35016 57152
rect 35080 57088 35096 57152
rect 35160 57088 35176 57152
rect 35240 57088 35248 57152
rect 34928 57087 35248 57088
rect 65648 57152 65968 57153
rect 65648 57088 65656 57152
rect 65720 57088 65736 57152
rect 65800 57088 65816 57152
rect 65880 57088 65896 57152
rect 65960 57088 65968 57152
rect 65648 57087 65968 57088
rect 19568 56608 19888 56609
rect 19568 56544 19576 56608
rect 19640 56544 19656 56608
rect 19720 56544 19736 56608
rect 19800 56544 19816 56608
rect 19880 56544 19888 56608
rect 19568 56543 19888 56544
rect 50288 56608 50608 56609
rect 50288 56544 50296 56608
rect 50360 56544 50376 56608
rect 50440 56544 50456 56608
rect 50520 56544 50536 56608
rect 50600 56544 50608 56608
rect 50288 56543 50608 56544
rect 4208 56064 4528 56065
rect 4208 56000 4216 56064
rect 4280 56000 4296 56064
rect 4360 56000 4376 56064
rect 4440 56000 4456 56064
rect 4520 56000 4528 56064
rect 4208 55999 4528 56000
rect 34928 56064 35248 56065
rect 34928 56000 34936 56064
rect 35000 56000 35016 56064
rect 35080 56000 35096 56064
rect 35160 56000 35176 56064
rect 35240 56000 35248 56064
rect 34928 55999 35248 56000
rect 65648 56064 65968 56065
rect 65648 56000 65656 56064
rect 65720 56000 65736 56064
rect 65800 56000 65816 56064
rect 65880 56000 65896 56064
rect 65960 56000 65968 56064
rect 65648 55999 65968 56000
rect 77845 55858 77911 55861
rect 79200 55858 80000 55888
rect 77845 55856 80000 55858
rect 77845 55800 77850 55856
rect 77906 55800 80000 55856
rect 77845 55798 80000 55800
rect 77845 55795 77911 55798
rect 79200 55768 80000 55798
rect 19568 55520 19888 55521
rect 19568 55456 19576 55520
rect 19640 55456 19656 55520
rect 19720 55456 19736 55520
rect 19800 55456 19816 55520
rect 19880 55456 19888 55520
rect 19568 55455 19888 55456
rect 50288 55520 50608 55521
rect 50288 55456 50296 55520
rect 50360 55456 50376 55520
rect 50440 55456 50456 55520
rect 50520 55456 50536 55520
rect 50600 55456 50608 55520
rect 50288 55455 50608 55456
rect 4208 54976 4528 54977
rect 4208 54912 4216 54976
rect 4280 54912 4296 54976
rect 4360 54912 4376 54976
rect 4440 54912 4456 54976
rect 4520 54912 4528 54976
rect 4208 54911 4528 54912
rect 34928 54976 35248 54977
rect 34928 54912 34936 54976
rect 35000 54912 35016 54976
rect 35080 54912 35096 54976
rect 35160 54912 35176 54976
rect 35240 54912 35248 54976
rect 34928 54911 35248 54912
rect 65648 54976 65968 54977
rect 65648 54912 65656 54976
rect 65720 54912 65736 54976
rect 65800 54912 65816 54976
rect 65880 54912 65896 54976
rect 65960 54912 65968 54976
rect 65648 54911 65968 54912
rect 0 54498 800 54528
rect 1485 54498 1551 54501
rect 0 54496 1551 54498
rect 0 54440 1490 54496
rect 1546 54440 1551 54496
rect 0 54438 1551 54440
rect 0 54408 800 54438
rect 1485 54435 1551 54438
rect 19568 54432 19888 54433
rect 19568 54368 19576 54432
rect 19640 54368 19656 54432
rect 19720 54368 19736 54432
rect 19800 54368 19816 54432
rect 19880 54368 19888 54432
rect 19568 54367 19888 54368
rect 50288 54432 50608 54433
rect 50288 54368 50296 54432
rect 50360 54368 50376 54432
rect 50440 54368 50456 54432
rect 50520 54368 50536 54432
rect 50600 54368 50608 54432
rect 50288 54367 50608 54368
rect 4208 53888 4528 53889
rect 4208 53824 4216 53888
rect 4280 53824 4296 53888
rect 4360 53824 4376 53888
rect 4440 53824 4456 53888
rect 4520 53824 4528 53888
rect 4208 53823 4528 53824
rect 34928 53888 35248 53889
rect 34928 53824 34936 53888
rect 35000 53824 35016 53888
rect 35080 53824 35096 53888
rect 35160 53824 35176 53888
rect 35240 53824 35248 53888
rect 34928 53823 35248 53824
rect 65648 53888 65968 53889
rect 65648 53824 65656 53888
rect 65720 53824 65736 53888
rect 65800 53824 65816 53888
rect 65880 53824 65896 53888
rect 65960 53824 65968 53888
rect 65648 53823 65968 53824
rect 19568 53344 19888 53345
rect 19568 53280 19576 53344
rect 19640 53280 19656 53344
rect 19720 53280 19736 53344
rect 19800 53280 19816 53344
rect 19880 53280 19888 53344
rect 19568 53279 19888 53280
rect 50288 53344 50608 53345
rect 50288 53280 50296 53344
rect 50360 53280 50376 53344
rect 50440 53280 50456 53344
rect 50520 53280 50536 53344
rect 50600 53280 50608 53344
rect 50288 53279 50608 53280
rect 4208 52800 4528 52801
rect 4208 52736 4216 52800
rect 4280 52736 4296 52800
rect 4360 52736 4376 52800
rect 4440 52736 4456 52800
rect 4520 52736 4528 52800
rect 4208 52735 4528 52736
rect 34928 52800 35248 52801
rect 34928 52736 34936 52800
rect 35000 52736 35016 52800
rect 35080 52736 35096 52800
rect 35160 52736 35176 52800
rect 35240 52736 35248 52800
rect 34928 52735 35248 52736
rect 65648 52800 65968 52801
rect 65648 52736 65656 52800
rect 65720 52736 65736 52800
rect 65800 52736 65816 52800
rect 65880 52736 65896 52800
rect 65960 52736 65968 52800
rect 65648 52735 65968 52736
rect 19568 52256 19888 52257
rect 19568 52192 19576 52256
rect 19640 52192 19656 52256
rect 19720 52192 19736 52256
rect 19800 52192 19816 52256
rect 19880 52192 19888 52256
rect 19568 52191 19888 52192
rect 50288 52256 50608 52257
rect 50288 52192 50296 52256
rect 50360 52192 50376 52256
rect 50440 52192 50456 52256
rect 50520 52192 50536 52256
rect 50600 52192 50608 52256
rect 50288 52191 50608 52192
rect 77845 51778 77911 51781
rect 79200 51778 80000 51808
rect 77845 51776 80000 51778
rect 77845 51720 77850 51776
rect 77906 51720 80000 51776
rect 77845 51718 80000 51720
rect 77845 51715 77911 51718
rect 4208 51712 4528 51713
rect 4208 51648 4216 51712
rect 4280 51648 4296 51712
rect 4360 51648 4376 51712
rect 4440 51648 4456 51712
rect 4520 51648 4528 51712
rect 4208 51647 4528 51648
rect 34928 51712 35248 51713
rect 34928 51648 34936 51712
rect 35000 51648 35016 51712
rect 35080 51648 35096 51712
rect 35160 51648 35176 51712
rect 35240 51648 35248 51712
rect 34928 51647 35248 51648
rect 65648 51712 65968 51713
rect 65648 51648 65656 51712
rect 65720 51648 65736 51712
rect 65800 51648 65816 51712
rect 65880 51648 65896 51712
rect 65960 51648 65968 51712
rect 79200 51688 80000 51718
rect 65648 51647 65968 51648
rect 19568 51168 19888 51169
rect 19568 51104 19576 51168
rect 19640 51104 19656 51168
rect 19720 51104 19736 51168
rect 19800 51104 19816 51168
rect 19880 51104 19888 51168
rect 19568 51103 19888 51104
rect 50288 51168 50608 51169
rect 50288 51104 50296 51168
rect 50360 51104 50376 51168
rect 50440 51104 50456 51168
rect 50520 51104 50536 51168
rect 50600 51104 50608 51168
rect 50288 51103 50608 51104
rect 4208 50624 4528 50625
rect 4208 50560 4216 50624
rect 4280 50560 4296 50624
rect 4360 50560 4376 50624
rect 4440 50560 4456 50624
rect 4520 50560 4528 50624
rect 4208 50559 4528 50560
rect 34928 50624 35248 50625
rect 34928 50560 34936 50624
rect 35000 50560 35016 50624
rect 35080 50560 35096 50624
rect 35160 50560 35176 50624
rect 35240 50560 35248 50624
rect 34928 50559 35248 50560
rect 65648 50624 65968 50625
rect 65648 50560 65656 50624
rect 65720 50560 65736 50624
rect 65800 50560 65816 50624
rect 65880 50560 65896 50624
rect 65960 50560 65968 50624
rect 65648 50559 65968 50560
rect 0 50418 800 50448
rect 1485 50418 1551 50421
rect 0 50416 1551 50418
rect 0 50360 1490 50416
rect 1546 50360 1551 50416
rect 0 50358 1551 50360
rect 0 50328 800 50358
rect 1485 50355 1551 50358
rect 19568 50080 19888 50081
rect 19568 50016 19576 50080
rect 19640 50016 19656 50080
rect 19720 50016 19736 50080
rect 19800 50016 19816 50080
rect 19880 50016 19888 50080
rect 19568 50015 19888 50016
rect 50288 50080 50608 50081
rect 50288 50016 50296 50080
rect 50360 50016 50376 50080
rect 50440 50016 50456 50080
rect 50520 50016 50536 50080
rect 50600 50016 50608 50080
rect 50288 50015 50608 50016
rect 4208 49536 4528 49537
rect 4208 49472 4216 49536
rect 4280 49472 4296 49536
rect 4360 49472 4376 49536
rect 4440 49472 4456 49536
rect 4520 49472 4528 49536
rect 4208 49471 4528 49472
rect 34928 49536 35248 49537
rect 34928 49472 34936 49536
rect 35000 49472 35016 49536
rect 35080 49472 35096 49536
rect 35160 49472 35176 49536
rect 35240 49472 35248 49536
rect 34928 49471 35248 49472
rect 65648 49536 65968 49537
rect 65648 49472 65656 49536
rect 65720 49472 65736 49536
rect 65800 49472 65816 49536
rect 65880 49472 65896 49536
rect 65960 49472 65968 49536
rect 65648 49471 65968 49472
rect 19568 48992 19888 48993
rect 19568 48928 19576 48992
rect 19640 48928 19656 48992
rect 19720 48928 19736 48992
rect 19800 48928 19816 48992
rect 19880 48928 19888 48992
rect 19568 48927 19888 48928
rect 50288 48992 50608 48993
rect 50288 48928 50296 48992
rect 50360 48928 50376 48992
rect 50440 48928 50456 48992
rect 50520 48928 50536 48992
rect 50600 48928 50608 48992
rect 50288 48927 50608 48928
rect 4208 48448 4528 48449
rect 4208 48384 4216 48448
rect 4280 48384 4296 48448
rect 4360 48384 4376 48448
rect 4440 48384 4456 48448
rect 4520 48384 4528 48448
rect 4208 48383 4528 48384
rect 34928 48448 35248 48449
rect 34928 48384 34936 48448
rect 35000 48384 35016 48448
rect 35080 48384 35096 48448
rect 35160 48384 35176 48448
rect 35240 48384 35248 48448
rect 34928 48383 35248 48384
rect 65648 48448 65968 48449
rect 65648 48384 65656 48448
rect 65720 48384 65736 48448
rect 65800 48384 65816 48448
rect 65880 48384 65896 48448
rect 65960 48384 65968 48448
rect 65648 48383 65968 48384
rect 19568 47904 19888 47905
rect 19568 47840 19576 47904
rect 19640 47840 19656 47904
rect 19720 47840 19736 47904
rect 19800 47840 19816 47904
rect 19880 47840 19888 47904
rect 19568 47839 19888 47840
rect 50288 47904 50608 47905
rect 50288 47840 50296 47904
rect 50360 47840 50376 47904
rect 50440 47840 50456 47904
rect 50520 47840 50536 47904
rect 50600 47840 50608 47904
rect 50288 47839 50608 47840
rect 75821 47698 75887 47701
rect 79200 47698 80000 47728
rect 75821 47696 80000 47698
rect 75821 47640 75826 47696
rect 75882 47640 80000 47696
rect 75821 47638 80000 47640
rect 75821 47635 75887 47638
rect 79200 47608 80000 47638
rect 4208 47360 4528 47361
rect 4208 47296 4216 47360
rect 4280 47296 4296 47360
rect 4360 47296 4376 47360
rect 4440 47296 4456 47360
rect 4520 47296 4528 47360
rect 4208 47295 4528 47296
rect 34928 47360 35248 47361
rect 34928 47296 34936 47360
rect 35000 47296 35016 47360
rect 35080 47296 35096 47360
rect 35160 47296 35176 47360
rect 35240 47296 35248 47360
rect 34928 47295 35248 47296
rect 65648 47360 65968 47361
rect 65648 47296 65656 47360
rect 65720 47296 65736 47360
rect 65800 47296 65816 47360
rect 65880 47296 65896 47360
rect 65960 47296 65968 47360
rect 65648 47295 65968 47296
rect 0 47018 800 47048
rect 1577 47018 1643 47021
rect 0 47016 1643 47018
rect 0 46960 1582 47016
rect 1638 46960 1643 47016
rect 0 46958 1643 46960
rect 0 46928 800 46958
rect 1577 46955 1643 46958
rect 19568 46816 19888 46817
rect 19568 46752 19576 46816
rect 19640 46752 19656 46816
rect 19720 46752 19736 46816
rect 19800 46752 19816 46816
rect 19880 46752 19888 46816
rect 19568 46751 19888 46752
rect 50288 46816 50608 46817
rect 50288 46752 50296 46816
rect 50360 46752 50376 46816
rect 50440 46752 50456 46816
rect 50520 46752 50536 46816
rect 50600 46752 50608 46816
rect 50288 46751 50608 46752
rect 4208 46272 4528 46273
rect 4208 46208 4216 46272
rect 4280 46208 4296 46272
rect 4360 46208 4376 46272
rect 4440 46208 4456 46272
rect 4520 46208 4528 46272
rect 4208 46207 4528 46208
rect 34928 46272 35248 46273
rect 34928 46208 34936 46272
rect 35000 46208 35016 46272
rect 35080 46208 35096 46272
rect 35160 46208 35176 46272
rect 35240 46208 35248 46272
rect 34928 46207 35248 46208
rect 65648 46272 65968 46273
rect 65648 46208 65656 46272
rect 65720 46208 65736 46272
rect 65800 46208 65816 46272
rect 65880 46208 65896 46272
rect 65960 46208 65968 46272
rect 65648 46207 65968 46208
rect 19568 45728 19888 45729
rect 19568 45664 19576 45728
rect 19640 45664 19656 45728
rect 19720 45664 19736 45728
rect 19800 45664 19816 45728
rect 19880 45664 19888 45728
rect 19568 45663 19888 45664
rect 50288 45728 50608 45729
rect 50288 45664 50296 45728
rect 50360 45664 50376 45728
rect 50440 45664 50456 45728
rect 50520 45664 50536 45728
rect 50600 45664 50608 45728
rect 50288 45663 50608 45664
rect 4208 45184 4528 45185
rect 4208 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4528 45184
rect 4208 45119 4528 45120
rect 34928 45184 35248 45185
rect 34928 45120 34936 45184
rect 35000 45120 35016 45184
rect 35080 45120 35096 45184
rect 35160 45120 35176 45184
rect 35240 45120 35248 45184
rect 34928 45119 35248 45120
rect 65648 45184 65968 45185
rect 65648 45120 65656 45184
rect 65720 45120 65736 45184
rect 65800 45120 65816 45184
rect 65880 45120 65896 45184
rect 65960 45120 65968 45184
rect 65648 45119 65968 45120
rect 19568 44640 19888 44641
rect 19568 44576 19576 44640
rect 19640 44576 19656 44640
rect 19720 44576 19736 44640
rect 19800 44576 19816 44640
rect 19880 44576 19888 44640
rect 19568 44575 19888 44576
rect 50288 44640 50608 44641
rect 50288 44576 50296 44640
rect 50360 44576 50376 44640
rect 50440 44576 50456 44640
rect 50520 44576 50536 44640
rect 50600 44576 50608 44640
rect 50288 44575 50608 44576
rect 4208 44096 4528 44097
rect 4208 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4528 44096
rect 4208 44031 4528 44032
rect 34928 44096 35248 44097
rect 34928 44032 34936 44096
rect 35000 44032 35016 44096
rect 35080 44032 35096 44096
rect 35160 44032 35176 44096
rect 35240 44032 35248 44096
rect 34928 44031 35248 44032
rect 65648 44096 65968 44097
rect 65648 44032 65656 44096
rect 65720 44032 65736 44096
rect 65800 44032 65816 44096
rect 65880 44032 65896 44096
rect 65960 44032 65968 44096
rect 65648 44031 65968 44032
rect 78029 43618 78095 43621
rect 79200 43618 80000 43648
rect 78029 43616 80000 43618
rect 78029 43560 78034 43616
rect 78090 43560 80000 43616
rect 78029 43558 80000 43560
rect 78029 43555 78095 43558
rect 19568 43552 19888 43553
rect 19568 43488 19576 43552
rect 19640 43488 19656 43552
rect 19720 43488 19736 43552
rect 19800 43488 19816 43552
rect 19880 43488 19888 43552
rect 19568 43487 19888 43488
rect 50288 43552 50608 43553
rect 50288 43488 50296 43552
rect 50360 43488 50376 43552
rect 50440 43488 50456 43552
rect 50520 43488 50536 43552
rect 50600 43488 50608 43552
rect 79200 43528 80000 43558
rect 50288 43487 50608 43488
rect 4208 43008 4528 43009
rect 0 42938 800 42968
rect 4208 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4528 43008
rect 4208 42943 4528 42944
rect 34928 43008 35248 43009
rect 34928 42944 34936 43008
rect 35000 42944 35016 43008
rect 35080 42944 35096 43008
rect 35160 42944 35176 43008
rect 35240 42944 35248 43008
rect 34928 42943 35248 42944
rect 65648 43008 65968 43009
rect 65648 42944 65656 43008
rect 65720 42944 65736 43008
rect 65800 42944 65816 43008
rect 65880 42944 65896 43008
rect 65960 42944 65968 43008
rect 65648 42943 65968 42944
rect 1853 42938 1919 42941
rect 0 42936 1919 42938
rect 0 42880 1858 42936
rect 1914 42880 1919 42936
rect 0 42878 1919 42880
rect 0 42848 800 42878
rect 1853 42875 1919 42878
rect 19568 42464 19888 42465
rect 19568 42400 19576 42464
rect 19640 42400 19656 42464
rect 19720 42400 19736 42464
rect 19800 42400 19816 42464
rect 19880 42400 19888 42464
rect 19568 42399 19888 42400
rect 50288 42464 50608 42465
rect 50288 42400 50296 42464
rect 50360 42400 50376 42464
rect 50440 42400 50456 42464
rect 50520 42400 50536 42464
rect 50600 42400 50608 42464
rect 50288 42399 50608 42400
rect 4208 41920 4528 41921
rect 4208 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4528 41920
rect 4208 41855 4528 41856
rect 34928 41920 35248 41921
rect 34928 41856 34936 41920
rect 35000 41856 35016 41920
rect 35080 41856 35096 41920
rect 35160 41856 35176 41920
rect 35240 41856 35248 41920
rect 34928 41855 35248 41856
rect 65648 41920 65968 41921
rect 65648 41856 65656 41920
rect 65720 41856 65736 41920
rect 65800 41856 65816 41920
rect 65880 41856 65896 41920
rect 65960 41856 65968 41920
rect 65648 41855 65968 41856
rect 19568 41376 19888 41377
rect 19568 41312 19576 41376
rect 19640 41312 19656 41376
rect 19720 41312 19736 41376
rect 19800 41312 19816 41376
rect 19880 41312 19888 41376
rect 19568 41311 19888 41312
rect 50288 41376 50608 41377
rect 50288 41312 50296 41376
rect 50360 41312 50376 41376
rect 50440 41312 50456 41376
rect 50520 41312 50536 41376
rect 50600 41312 50608 41376
rect 50288 41311 50608 41312
rect 4208 40832 4528 40833
rect 4208 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4528 40832
rect 4208 40767 4528 40768
rect 34928 40832 35248 40833
rect 34928 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35248 40832
rect 34928 40767 35248 40768
rect 65648 40832 65968 40833
rect 65648 40768 65656 40832
rect 65720 40768 65736 40832
rect 65800 40768 65816 40832
rect 65880 40768 65896 40832
rect 65960 40768 65968 40832
rect 65648 40767 65968 40768
rect 19568 40288 19888 40289
rect 19568 40224 19576 40288
rect 19640 40224 19656 40288
rect 19720 40224 19736 40288
rect 19800 40224 19816 40288
rect 19880 40224 19888 40288
rect 19568 40223 19888 40224
rect 50288 40288 50608 40289
rect 50288 40224 50296 40288
rect 50360 40224 50376 40288
rect 50440 40224 50456 40288
rect 50520 40224 50536 40288
rect 50600 40224 50608 40288
rect 50288 40223 50608 40224
rect 78029 40218 78095 40221
rect 79200 40218 80000 40248
rect 78029 40216 80000 40218
rect 78029 40160 78034 40216
rect 78090 40160 80000 40216
rect 78029 40158 80000 40160
rect 78029 40155 78095 40158
rect 79200 40128 80000 40158
rect 4208 39744 4528 39745
rect 4208 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4528 39744
rect 4208 39679 4528 39680
rect 34928 39744 35248 39745
rect 34928 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35248 39744
rect 34928 39679 35248 39680
rect 65648 39744 65968 39745
rect 65648 39680 65656 39744
rect 65720 39680 65736 39744
rect 65800 39680 65816 39744
rect 65880 39680 65896 39744
rect 65960 39680 65968 39744
rect 65648 39679 65968 39680
rect 19568 39200 19888 39201
rect 19568 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19888 39200
rect 19568 39135 19888 39136
rect 50288 39200 50608 39201
rect 50288 39136 50296 39200
rect 50360 39136 50376 39200
rect 50440 39136 50456 39200
rect 50520 39136 50536 39200
rect 50600 39136 50608 39200
rect 50288 39135 50608 39136
rect 0 38858 800 38888
rect 1853 38858 1919 38861
rect 0 38856 1919 38858
rect 0 38800 1858 38856
rect 1914 38800 1919 38856
rect 0 38798 1919 38800
rect 0 38768 800 38798
rect 1853 38795 1919 38798
rect 4208 38656 4528 38657
rect 4208 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4528 38656
rect 4208 38591 4528 38592
rect 34928 38656 35248 38657
rect 34928 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35248 38656
rect 34928 38591 35248 38592
rect 65648 38656 65968 38657
rect 65648 38592 65656 38656
rect 65720 38592 65736 38656
rect 65800 38592 65816 38656
rect 65880 38592 65896 38656
rect 65960 38592 65968 38656
rect 65648 38591 65968 38592
rect 19568 38112 19888 38113
rect 19568 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19888 38112
rect 19568 38047 19888 38048
rect 50288 38112 50608 38113
rect 50288 38048 50296 38112
rect 50360 38048 50376 38112
rect 50440 38048 50456 38112
rect 50520 38048 50536 38112
rect 50600 38048 50608 38112
rect 50288 38047 50608 38048
rect 4208 37568 4528 37569
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 37503 4528 37504
rect 34928 37568 35248 37569
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 37503 35248 37504
rect 65648 37568 65968 37569
rect 65648 37504 65656 37568
rect 65720 37504 65736 37568
rect 65800 37504 65816 37568
rect 65880 37504 65896 37568
rect 65960 37504 65968 37568
rect 65648 37503 65968 37504
rect 19568 37024 19888 37025
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 36959 19888 36960
rect 50288 37024 50608 37025
rect 50288 36960 50296 37024
rect 50360 36960 50376 37024
rect 50440 36960 50456 37024
rect 50520 36960 50536 37024
rect 50600 36960 50608 37024
rect 50288 36959 50608 36960
rect 4208 36480 4528 36481
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 36415 4528 36416
rect 34928 36480 35248 36481
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 36415 35248 36416
rect 65648 36480 65968 36481
rect 65648 36416 65656 36480
rect 65720 36416 65736 36480
rect 65800 36416 65816 36480
rect 65880 36416 65896 36480
rect 65960 36416 65968 36480
rect 65648 36415 65968 36416
rect 78029 36138 78095 36141
rect 79200 36138 80000 36168
rect 78029 36136 80000 36138
rect 78029 36080 78034 36136
rect 78090 36080 80000 36136
rect 78029 36078 80000 36080
rect 78029 36075 78095 36078
rect 79200 36048 80000 36078
rect 19568 35936 19888 35937
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 35871 19888 35872
rect 50288 35936 50608 35937
rect 50288 35872 50296 35936
rect 50360 35872 50376 35936
rect 50440 35872 50456 35936
rect 50520 35872 50536 35936
rect 50600 35872 50608 35936
rect 50288 35871 50608 35872
rect 4208 35392 4528 35393
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 35327 4528 35328
rect 34928 35392 35248 35393
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 35327 35248 35328
rect 65648 35392 65968 35393
rect 65648 35328 65656 35392
rect 65720 35328 65736 35392
rect 65800 35328 65816 35392
rect 65880 35328 65896 35392
rect 65960 35328 65968 35392
rect 65648 35327 65968 35328
rect 19568 34848 19888 34849
rect 0 34778 800 34808
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 34783 19888 34784
rect 50288 34848 50608 34849
rect 50288 34784 50296 34848
rect 50360 34784 50376 34848
rect 50440 34784 50456 34848
rect 50520 34784 50536 34848
rect 50600 34784 50608 34848
rect 50288 34783 50608 34784
rect 1577 34778 1643 34781
rect 0 34776 1643 34778
rect 0 34720 1582 34776
rect 1638 34720 1643 34776
rect 0 34718 1643 34720
rect 0 34688 800 34718
rect 1577 34715 1643 34718
rect 4208 34304 4528 34305
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 34239 4528 34240
rect 34928 34304 35248 34305
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 34239 35248 34240
rect 65648 34304 65968 34305
rect 65648 34240 65656 34304
rect 65720 34240 65736 34304
rect 65800 34240 65816 34304
rect 65880 34240 65896 34304
rect 65960 34240 65968 34304
rect 65648 34239 65968 34240
rect 19568 33760 19888 33761
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 33695 19888 33696
rect 50288 33760 50608 33761
rect 50288 33696 50296 33760
rect 50360 33696 50376 33760
rect 50440 33696 50456 33760
rect 50520 33696 50536 33760
rect 50600 33696 50608 33760
rect 50288 33695 50608 33696
rect 4208 33216 4528 33217
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 33151 4528 33152
rect 34928 33216 35248 33217
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 33151 35248 33152
rect 65648 33216 65968 33217
rect 65648 33152 65656 33216
rect 65720 33152 65736 33216
rect 65800 33152 65816 33216
rect 65880 33152 65896 33216
rect 65960 33152 65968 33216
rect 65648 33151 65968 33152
rect 19568 32672 19888 32673
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 32607 19888 32608
rect 50288 32672 50608 32673
rect 50288 32608 50296 32672
rect 50360 32608 50376 32672
rect 50440 32608 50456 32672
rect 50520 32608 50536 32672
rect 50600 32608 50608 32672
rect 50288 32607 50608 32608
rect 4208 32128 4528 32129
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 32063 4528 32064
rect 34928 32128 35248 32129
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 32063 35248 32064
rect 65648 32128 65968 32129
rect 65648 32064 65656 32128
rect 65720 32064 65736 32128
rect 65800 32064 65816 32128
rect 65880 32064 65896 32128
rect 65960 32064 65968 32128
rect 65648 32063 65968 32064
rect 77753 32058 77819 32061
rect 79200 32058 80000 32088
rect 77753 32056 80000 32058
rect 77753 32000 77758 32056
rect 77814 32000 80000 32056
rect 77753 31998 80000 32000
rect 77753 31995 77819 31998
rect 79200 31968 80000 31998
rect 19568 31584 19888 31585
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 31519 19888 31520
rect 50288 31584 50608 31585
rect 50288 31520 50296 31584
rect 50360 31520 50376 31584
rect 50440 31520 50456 31584
rect 50520 31520 50536 31584
rect 50600 31520 50608 31584
rect 50288 31519 50608 31520
rect 0 31378 800 31408
rect 1393 31378 1459 31381
rect 0 31376 1459 31378
rect 0 31320 1398 31376
rect 1454 31320 1459 31376
rect 0 31318 1459 31320
rect 0 31288 800 31318
rect 1393 31315 1459 31318
rect 4208 31040 4528 31041
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 30975 4528 30976
rect 34928 31040 35248 31041
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 30975 35248 30976
rect 65648 31040 65968 31041
rect 65648 30976 65656 31040
rect 65720 30976 65736 31040
rect 65800 30976 65816 31040
rect 65880 30976 65896 31040
rect 65960 30976 65968 31040
rect 65648 30975 65968 30976
rect 19568 30496 19888 30497
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 30431 19888 30432
rect 50288 30496 50608 30497
rect 50288 30432 50296 30496
rect 50360 30432 50376 30496
rect 50440 30432 50456 30496
rect 50520 30432 50536 30496
rect 50600 30432 50608 30496
rect 50288 30431 50608 30432
rect 4208 29952 4528 29953
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 29887 4528 29888
rect 34928 29952 35248 29953
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 29887 35248 29888
rect 65648 29952 65968 29953
rect 65648 29888 65656 29952
rect 65720 29888 65736 29952
rect 65800 29888 65816 29952
rect 65880 29888 65896 29952
rect 65960 29888 65968 29952
rect 65648 29887 65968 29888
rect 19568 29408 19888 29409
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 29343 19888 29344
rect 50288 29408 50608 29409
rect 50288 29344 50296 29408
rect 50360 29344 50376 29408
rect 50440 29344 50456 29408
rect 50520 29344 50536 29408
rect 50600 29344 50608 29408
rect 50288 29343 50608 29344
rect 4208 28864 4528 28865
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 28799 4528 28800
rect 34928 28864 35248 28865
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 28799 35248 28800
rect 65648 28864 65968 28865
rect 65648 28800 65656 28864
rect 65720 28800 65736 28864
rect 65800 28800 65816 28864
rect 65880 28800 65896 28864
rect 65960 28800 65968 28864
rect 65648 28799 65968 28800
rect 19568 28320 19888 28321
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 28255 19888 28256
rect 50288 28320 50608 28321
rect 50288 28256 50296 28320
rect 50360 28256 50376 28320
rect 50440 28256 50456 28320
rect 50520 28256 50536 28320
rect 50600 28256 50608 28320
rect 50288 28255 50608 28256
rect 77937 27978 78003 27981
rect 79200 27978 80000 28008
rect 77937 27976 80000 27978
rect 77937 27920 77942 27976
rect 77998 27920 80000 27976
rect 77937 27918 80000 27920
rect 77937 27915 78003 27918
rect 79200 27888 80000 27918
rect 4208 27776 4528 27777
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 27711 4528 27712
rect 34928 27776 35248 27777
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 27711 35248 27712
rect 65648 27776 65968 27777
rect 65648 27712 65656 27776
rect 65720 27712 65736 27776
rect 65800 27712 65816 27776
rect 65880 27712 65896 27776
rect 65960 27712 65968 27776
rect 65648 27711 65968 27712
rect 0 27298 800 27328
rect 1393 27298 1459 27301
rect 0 27296 1459 27298
rect 0 27240 1398 27296
rect 1454 27240 1459 27296
rect 0 27238 1459 27240
rect 0 27208 800 27238
rect 1393 27235 1459 27238
rect 19568 27232 19888 27233
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 27167 19888 27168
rect 50288 27232 50608 27233
rect 50288 27168 50296 27232
rect 50360 27168 50376 27232
rect 50440 27168 50456 27232
rect 50520 27168 50536 27232
rect 50600 27168 50608 27232
rect 50288 27167 50608 27168
rect 4208 26688 4528 26689
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 26623 4528 26624
rect 34928 26688 35248 26689
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 26623 35248 26624
rect 65648 26688 65968 26689
rect 65648 26624 65656 26688
rect 65720 26624 65736 26688
rect 65800 26624 65816 26688
rect 65880 26624 65896 26688
rect 65960 26624 65968 26688
rect 65648 26623 65968 26624
rect 19568 26144 19888 26145
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 26079 19888 26080
rect 50288 26144 50608 26145
rect 50288 26080 50296 26144
rect 50360 26080 50376 26144
rect 50440 26080 50456 26144
rect 50520 26080 50536 26144
rect 50600 26080 50608 26144
rect 50288 26079 50608 26080
rect 4208 25600 4528 25601
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 25535 4528 25536
rect 34928 25600 35248 25601
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 25535 35248 25536
rect 65648 25600 65968 25601
rect 65648 25536 65656 25600
rect 65720 25536 65736 25600
rect 65800 25536 65816 25600
rect 65880 25536 65896 25600
rect 65960 25536 65968 25600
rect 65648 25535 65968 25536
rect 19568 25056 19888 25057
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 24991 19888 24992
rect 50288 25056 50608 25057
rect 50288 24992 50296 25056
rect 50360 24992 50376 25056
rect 50440 24992 50456 25056
rect 50520 24992 50536 25056
rect 50600 24992 50608 25056
rect 50288 24991 50608 24992
rect 77845 24578 77911 24581
rect 79200 24578 80000 24608
rect 77845 24576 80000 24578
rect 77845 24520 77850 24576
rect 77906 24520 80000 24576
rect 77845 24518 80000 24520
rect 77845 24515 77911 24518
rect 4208 24512 4528 24513
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 24447 4528 24448
rect 34928 24512 35248 24513
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 24447 35248 24448
rect 65648 24512 65968 24513
rect 65648 24448 65656 24512
rect 65720 24448 65736 24512
rect 65800 24448 65816 24512
rect 65880 24448 65896 24512
rect 65960 24448 65968 24512
rect 79200 24488 80000 24518
rect 65648 24447 65968 24448
rect 19568 23968 19888 23969
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 23903 19888 23904
rect 50288 23968 50608 23969
rect 50288 23904 50296 23968
rect 50360 23904 50376 23968
rect 50440 23904 50456 23968
rect 50520 23904 50536 23968
rect 50600 23904 50608 23968
rect 50288 23903 50608 23904
rect 4208 23424 4528 23425
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 23359 4528 23360
rect 34928 23424 35248 23425
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 23359 35248 23360
rect 65648 23424 65968 23425
rect 65648 23360 65656 23424
rect 65720 23360 65736 23424
rect 65800 23360 65816 23424
rect 65880 23360 65896 23424
rect 65960 23360 65968 23424
rect 65648 23359 65968 23360
rect 0 23218 800 23248
rect 1393 23218 1459 23221
rect 0 23216 1459 23218
rect 0 23160 1398 23216
rect 1454 23160 1459 23216
rect 0 23158 1459 23160
rect 0 23128 800 23158
rect 1393 23155 1459 23158
rect 19568 22880 19888 22881
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 22815 19888 22816
rect 50288 22880 50608 22881
rect 50288 22816 50296 22880
rect 50360 22816 50376 22880
rect 50440 22816 50456 22880
rect 50520 22816 50536 22880
rect 50600 22816 50608 22880
rect 50288 22815 50608 22816
rect 4208 22336 4528 22337
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 22271 4528 22272
rect 34928 22336 35248 22337
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 22271 35248 22272
rect 65648 22336 65968 22337
rect 65648 22272 65656 22336
rect 65720 22272 65736 22336
rect 65800 22272 65816 22336
rect 65880 22272 65896 22336
rect 65960 22272 65968 22336
rect 65648 22271 65968 22272
rect 19568 21792 19888 21793
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 21727 19888 21728
rect 50288 21792 50608 21793
rect 50288 21728 50296 21792
rect 50360 21728 50376 21792
rect 50440 21728 50456 21792
rect 50520 21728 50536 21792
rect 50600 21728 50608 21792
rect 50288 21727 50608 21728
rect 4208 21248 4528 21249
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 21183 4528 21184
rect 34928 21248 35248 21249
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 21183 35248 21184
rect 65648 21248 65968 21249
rect 65648 21184 65656 21248
rect 65720 21184 65736 21248
rect 65800 21184 65816 21248
rect 65880 21184 65896 21248
rect 65960 21184 65968 21248
rect 65648 21183 65968 21184
rect 19568 20704 19888 20705
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 20639 19888 20640
rect 50288 20704 50608 20705
rect 50288 20640 50296 20704
rect 50360 20640 50376 20704
rect 50440 20640 50456 20704
rect 50520 20640 50536 20704
rect 50600 20640 50608 20704
rect 50288 20639 50608 20640
rect 78029 20498 78095 20501
rect 79200 20498 80000 20528
rect 78029 20496 80000 20498
rect 78029 20440 78034 20496
rect 78090 20440 80000 20496
rect 78029 20438 80000 20440
rect 78029 20435 78095 20438
rect 79200 20408 80000 20438
rect 4208 20160 4528 20161
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 20095 4528 20096
rect 34928 20160 35248 20161
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 20095 35248 20096
rect 65648 20160 65968 20161
rect 65648 20096 65656 20160
rect 65720 20096 65736 20160
rect 65800 20096 65816 20160
rect 65880 20096 65896 20160
rect 65960 20096 65968 20160
rect 65648 20095 65968 20096
rect 19568 19616 19888 19617
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 19551 19888 19552
rect 50288 19616 50608 19617
rect 50288 19552 50296 19616
rect 50360 19552 50376 19616
rect 50440 19552 50456 19616
rect 50520 19552 50536 19616
rect 50600 19552 50608 19616
rect 50288 19551 50608 19552
rect 0 19138 800 19168
rect 1577 19138 1643 19141
rect 0 19136 1643 19138
rect 0 19080 1582 19136
rect 1638 19080 1643 19136
rect 0 19078 1643 19080
rect 0 19048 800 19078
rect 1577 19075 1643 19078
rect 4208 19072 4528 19073
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 19007 4528 19008
rect 34928 19072 35248 19073
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 19007 35248 19008
rect 65648 19072 65968 19073
rect 65648 19008 65656 19072
rect 65720 19008 65736 19072
rect 65800 19008 65816 19072
rect 65880 19008 65896 19072
rect 65960 19008 65968 19072
rect 65648 19007 65968 19008
rect 19568 18528 19888 18529
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 18463 19888 18464
rect 50288 18528 50608 18529
rect 50288 18464 50296 18528
rect 50360 18464 50376 18528
rect 50440 18464 50456 18528
rect 50520 18464 50536 18528
rect 50600 18464 50608 18528
rect 50288 18463 50608 18464
rect 4208 17984 4528 17985
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 17919 4528 17920
rect 34928 17984 35248 17985
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 17919 35248 17920
rect 65648 17984 65968 17985
rect 65648 17920 65656 17984
rect 65720 17920 65736 17984
rect 65800 17920 65816 17984
rect 65880 17920 65896 17984
rect 65960 17920 65968 17984
rect 65648 17919 65968 17920
rect 19568 17440 19888 17441
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 17375 19888 17376
rect 50288 17440 50608 17441
rect 50288 17376 50296 17440
rect 50360 17376 50376 17440
rect 50440 17376 50456 17440
rect 50520 17376 50536 17440
rect 50600 17376 50608 17440
rect 50288 17375 50608 17376
rect 4208 16896 4528 16897
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 16831 4528 16832
rect 34928 16896 35248 16897
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 16831 35248 16832
rect 65648 16896 65968 16897
rect 65648 16832 65656 16896
rect 65720 16832 65736 16896
rect 65800 16832 65816 16896
rect 65880 16832 65896 16896
rect 65960 16832 65968 16896
rect 65648 16831 65968 16832
rect 78029 16418 78095 16421
rect 79200 16418 80000 16448
rect 78029 16416 80000 16418
rect 78029 16360 78034 16416
rect 78090 16360 80000 16416
rect 78029 16358 80000 16360
rect 78029 16355 78095 16358
rect 19568 16352 19888 16353
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 16287 19888 16288
rect 50288 16352 50608 16353
rect 50288 16288 50296 16352
rect 50360 16288 50376 16352
rect 50440 16288 50456 16352
rect 50520 16288 50536 16352
rect 50600 16288 50608 16352
rect 79200 16328 80000 16358
rect 50288 16287 50608 16288
rect 4208 15808 4528 15809
rect 0 15738 800 15768
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 15743 4528 15744
rect 34928 15808 35248 15809
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 15743 35248 15744
rect 65648 15808 65968 15809
rect 65648 15744 65656 15808
rect 65720 15744 65736 15808
rect 65800 15744 65816 15808
rect 65880 15744 65896 15808
rect 65960 15744 65968 15808
rect 65648 15743 65968 15744
rect 1485 15738 1551 15741
rect 0 15736 1551 15738
rect 0 15680 1490 15736
rect 1546 15680 1551 15736
rect 0 15678 1551 15680
rect 0 15648 800 15678
rect 1485 15675 1551 15678
rect 19568 15264 19888 15265
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 15199 19888 15200
rect 50288 15264 50608 15265
rect 50288 15200 50296 15264
rect 50360 15200 50376 15264
rect 50440 15200 50456 15264
rect 50520 15200 50536 15264
rect 50600 15200 50608 15264
rect 50288 15199 50608 15200
rect 4208 14720 4528 14721
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 14655 4528 14656
rect 34928 14720 35248 14721
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 14655 35248 14656
rect 65648 14720 65968 14721
rect 65648 14656 65656 14720
rect 65720 14656 65736 14720
rect 65800 14656 65816 14720
rect 65880 14656 65896 14720
rect 65960 14656 65968 14720
rect 65648 14655 65968 14656
rect 19568 14176 19888 14177
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 14111 19888 14112
rect 50288 14176 50608 14177
rect 50288 14112 50296 14176
rect 50360 14112 50376 14176
rect 50440 14112 50456 14176
rect 50520 14112 50536 14176
rect 50600 14112 50608 14176
rect 50288 14111 50608 14112
rect 4208 13632 4528 13633
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 13567 4528 13568
rect 34928 13632 35248 13633
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 13567 35248 13568
rect 65648 13632 65968 13633
rect 65648 13568 65656 13632
rect 65720 13568 65736 13632
rect 65800 13568 65816 13632
rect 65880 13568 65896 13632
rect 65960 13568 65968 13632
rect 65648 13567 65968 13568
rect 19568 13088 19888 13089
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 13023 19888 13024
rect 50288 13088 50608 13089
rect 50288 13024 50296 13088
rect 50360 13024 50376 13088
rect 50440 13024 50456 13088
rect 50520 13024 50536 13088
rect 50600 13024 50608 13088
rect 50288 13023 50608 13024
rect 4208 12544 4528 12545
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 12479 4528 12480
rect 34928 12544 35248 12545
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 12479 35248 12480
rect 65648 12544 65968 12545
rect 65648 12480 65656 12544
rect 65720 12480 65736 12544
rect 65800 12480 65816 12544
rect 65880 12480 65896 12544
rect 65960 12480 65968 12544
rect 65648 12479 65968 12480
rect 77201 12338 77267 12341
rect 79200 12338 80000 12368
rect 77201 12336 80000 12338
rect 77201 12280 77206 12336
rect 77262 12280 80000 12336
rect 77201 12278 80000 12280
rect 77201 12275 77267 12278
rect 79200 12248 80000 12278
rect 19568 12000 19888 12001
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 11935 19888 11936
rect 50288 12000 50608 12001
rect 50288 11936 50296 12000
rect 50360 11936 50376 12000
rect 50440 11936 50456 12000
rect 50520 11936 50536 12000
rect 50600 11936 50608 12000
rect 50288 11935 50608 11936
rect 0 11658 800 11688
rect 1393 11658 1459 11661
rect 0 11656 1459 11658
rect 0 11600 1398 11656
rect 1454 11600 1459 11656
rect 0 11598 1459 11600
rect 0 11568 800 11598
rect 1393 11595 1459 11598
rect 4208 11456 4528 11457
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 11391 4528 11392
rect 34928 11456 35248 11457
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 11391 35248 11392
rect 65648 11456 65968 11457
rect 65648 11392 65656 11456
rect 65720 11392 65736 11456
rect 65800 11392 65816 11456
rect 65880 11392 65896 11456
rect 65960 11392 65968 11456
rect 65648 11391 65968 11392
rect 19568 10912 19888 10913
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 10847 19888 10848
rect 50288 10912 50608 10913
rect 50288 10848 50296 10912
rect 50360 10848 50376 10912
rect 50440 10848 50456 10912
rect 50520 10848 50536 10912
rect 50600 10848 50608 10912
rect 50288 10847 50608 10848
rect 4208 10368 4528 10369
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 10303 4528 10304
rect 34928 10368 35248 10369
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 10303 35248 10304
rect 65648 10368 65968 10369
rect 65648 10304 65656 10368
rect 65720 10304 65736 10368
rect 65800 10304 65816 10368
rect 65880 10304 65896 10368
rect 65960 10304 65968 10368
rect 65648 10303 65968 10304
rect 19568 9824 19888 9825
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 9759 19888 9760
rect 50288 9824 50608 9825
rect 50288 9760 50296 9824
rect 50360 9760 50376 9824
rect 50440 9760 50456 9824
rect 50520 9760 50536 9824
rect 50600 9760 50608 9824
rect 50288 9759 50608 9760
rect 4208 9280 4528 9281
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 9215 4528 9216
rect 34928 9280 35248 9281
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 9215 35248 9216
rect 65648 9280 65968 9281
rect 65648 9216 65656 9280
rect 65720 9216 65736 9280
rect 65800 9216 65816 9280
rect 65880 9216 65896 9280
rect 65960 9216 65968 9280
rect 65648 9215 65968 9216
rect 78029 8938 78095 8941
rect 79200 8938 80000 8968
rect 78029 8936 80000 8938
rect 78029 8880 78034 8936
rect 78090 8880 80000 8936
rect 78029 8878 80000 8880
rect 78029 8875 78095 8878
rect 79200 8848 80000 8878
rect 19568 8736 19888 8737
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 8671 19888 8672
rect 50288 8736 50608 8737
rect 50288 8672 50296 8736
rect 50360 8672 50376 8736
rect 50440 8672 50456 8736
rect 50520 8672 50536 8736
rect 50600 8672 50608 8736
rect 50288 8671 50608 8672
rect 4208 8192 4528 8193
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 8127 4528 8128
rect 34928 8192 35248 8193
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 8127 35248 8128
rect 65648 8192 65968 8193
rect 65648 8128 65656 8192
rect 65720 8128 65736 8192
rect 65800 8128 65816 8192
rect 65880 8128 65896 8192
rect 65960 8128 65968 8192
rect 65648 8127 65968 8128
rect 19568 7648 19888 7649
rect 0 7578 800 7608
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 7583 19888 7584
rect 50288 7648 50608 7649
rect 50288 7584 50296 7648
rect 50360 7584 50376 7648
rect 50440 7584 50456 7648
rect 50520 7584 50536 7648
rect 50600 7584 50608 7648
rect 50288 7583 50608 7584
rect 1577 7578 1643 7581
rect 0 7576 1643 7578
rect 0 7520 1582 7576
rect 1638 7520 1643 7576
rect 0 7518 1643 7520
rect 0 7488 800 7518
rect 1577 7515 1643 7518
rect 4208 7104 4528 7105
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 7039 4528 7040
rect 34928 7104 35248 7105
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 7039 35248 7040
rect 65648 7104 65968 7105
rect 65648 7040 65656 7104
rect 65720 7040 65736 7104
rect 65800 7040 65816 7104
rect 65880 7040 65896 7104
rect 65960 7040 65968 7104
rect 65648 7039 65968 7040
rect 19568 6560 19888 6561
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 6495 19888 6496
rect 50288 6560 50608 6561
rect 50288 6496 50296 6560
rect 50360 6496 50376 6560
rect 50440 6496 50456 6560
rect 50520 6496 50536 6560
rect 50600 6496 50608 6560
rect 50288 6495 50608 6496
rect 4208 6016 4528 6017
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 5951 4528 5952
rect 34928 6016 35248 6017
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 5951 35248 5952
rect 65648 6016 65968 6017
rect 65648 5952 65656 6016
rect 65720 5952 65736 6016
rect 65800 5952 65816 6016
rect 65880 5952 65896 6016
rect 65960 5952 65968 6016
rect 65648 5951 65968 5952
rect 19568 5472 19888 5473
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 5407 19888 5408
rect 50288 5472 50608 5473
rect 50288 5408 50296 5472
rect 50360 5408 50376 5472
rect 50440 5408 50456 5472
rect 50520 5408 50536 5472
rect 50600 5408 50608 5472
rect 50288 5407 50608 5408
rect 4208 4928 4528 4929
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 4863 4528 4864
rect 34928 4928 35248 4929
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 4863 35248 4864
rect 65648 4928 65968 4929
rect 65648 4864 65656 4928
rect 65720 4864 65736 4928
rect 65800 4864 65816 4928
rect 65880 4864 65896 4928
rect 65960 4864 65968 4928
rect 65648 4863 65968 4864
rect 77845 4858 77911 4861
rect 79200 4858 80000 4888
rect 77845 4856 80000 4858
rect 77845 4800 77850 4856
rect 77906 4800 80000 4856
rect 77845 4798 80000 4800
rect 77845 4795 77911 4798
rect 79200 4768 80000 4798
rect 19568 4384 19888 4385
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 4319 19888 4320
rect 50288 4384 50608 4385
rect 50288 4320 50296 4384
rect 50360 4320 50376 4384
rect 50440 4320 50456 4384
rect 50520 4320 50536 4384
rect 50600 4320 50608 4384
rect 50288 4319 50608 4320
rect 4208 3840 4528 3841
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 3775 4528 3776
rect 34928 3840 35248 3841
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 3775 35248 3776
rect 65648 3840 65968 3841
rect 65648 3776 65656 3840
rect 65720 3776 65736 3840
rect 65800 3776 65816 3840
rect 65880 3776 65896 3840
rect 65960 3776 65968 3840
rect 65648 3775 65968 3776
rect 0 3498 800 3528
rect 1393 3498 1459 3501
rect 0 3496 1459 3498
rect 0 3440 1398 3496
rect 1454 3440 1459 3496
rect 0 3438 1459 3440
rect 0 3408 800 3438
rect 1393 3435 1459 3438
rect 19568 3296 19888 3297
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19568 3231 19888 3232
rect 50288 3296 50608 3297
rect 50288 3232 50296 3296
rect 50360 3232 50376 3296
rect 50440 3232 50456 3296
rect 50520 3232 50536 3296
rect 50600 3232 50608 3296
rect 50288 3231 50608 3232
rect 4208 2752 4528 2753
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2687 4528 2688
rect 34928 2752 35248 2753
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2687 35248 2688
rect 65648 2752 65968 2753
rect 65648 2688 65656 2752
rect 65720 2688 65736 2752
rect 65800 2688 65816 2752
rect 65880 2688 65896 2752
rect 65960 2688 65968 2752
rect 65648 2687 65968 2688
rect 19568 2208 19888 2209
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2143 19888 2144
rect 50288 2208 50608 2209
rect 50288 2144 50296 2208
rect 50360 2144 50376 2208
rect 50440 2144 50456 2208
rect 50520 2144 50536 2208
rect 50600 2144 50608 2208
rect 50288 2143 50608 2144
rect 77661 778 77727 781
rect 79200 778 80000 808
rect 77661 776 80000 778
rect 77661 720 77666 776
rect 77722 720 80000 776
rect 77661 718 80000 720
rect 77661 715 77727 718
rect 79200 688 80000 718
<< via3 >>
rect 19576 117532 19640 117536
rect 19576 117476 19580 117532
rect 19580 117476 19636 117532
rect 19636 117476 19640 117532
rect 19576 117472 19640 117476
rect 19656 117532 19720 117536
rect 19656 117476 19660 117532
rect 19660 117476 19716 117532
rect 19716 117476 19720 117532
rect 19656 117472 19720 117476
rect 19736 117532 19800 117536
rect 19736 117476 19740 117532
rect 19740 117476 19796 117532
rect 19796 117476 19800 117532
rect 19736 117472 19800 117476
rect 19816 117532 19880 117536
rect 19816 117476 19820 117532
rect 19820 117476 19876 117532
rect 19876 117476 19880 117532
rect 19816 117472 19880 117476
rect 50296 117532 50360 117536
rect 50296 117476 50300 117532
rect 50300 117476 50356 117532
rect 50356 117476 50360 117532
rect 50296 117472 50360 117476
rect 50376 117532 50440 117536
rect 50376 117476 50380 117532
rect 50380 117476 50436 117532
rect 50436 117476 50440 117532
rect 50376 117472 50440 117476
rect 50456 117532 50520 117536
rect 50456 117476 50460 117532
rect 50460 117476 50516 117532
rect 50516 117476 50520 117532
rect 50456 117472 50520 117476
rect 50536 117532 50600 117536
rect 50536 117476 50540 117532
rect 50540 117476 50596 117532
rect 50596 117476 50600 117532
rect 50536 117472 50600 117476
rect 4216 116988 4280 116992
rect 4216 116932 4220 116988
rect 4220 116932 4276 116988
rect 4276 116932 4280 116988
rect 4216 116928 4280 116932
rect 4296 116988 4360 116992
rect 4296 116932 4300 116988
rect 4300 116932 4356 116988
rect 4356 116932 4360 116988
rect 4296 116928 4360 116932
rect 4376 116988 4440 116992
rect 4376 116932 4380 116988
rect 4380 116932 4436 116988
rect 4436 116932 4440 116988
rect 4376 116928 4440 116932
rect 4456 116988 4520 116992
rect 4456 116932 4460 116988
rect 4460 116932 4516 116988
rect 4516 116932 4520 116988
rect 4456 116928 4520 116932
rect 34936 116988 35000 116992
rect 34936 116932 34940 116988
rect 34940 116932 34996 116988
rect 34996 116932 35000 116988
rect 34936 116928 35000 116932
rect 35016 116988 35080 116992
rect 35016 116932 35020 116988
rect 35020 116932 35076 116988
rect 35076 116932 35080 116988
rect 35016 116928 35080 116932
rect 35096 116988 35160 116992
rect 35096 116932 35100 116988
rect 35100 116932 35156 116988
rect 35156 116932 35160 116988
rect 35096 116928 35160 116932
rect 35176 116988 35240 116992
rect 35176 116932 35180 116988
rect 35180 116932 35236 116988
rect 35236 116932 35240 116988
rect 35176 116928 35240 116932
rect 65656 116988 65720 116992
rect 65656 116932 65660 116988
rect 65660 116932 65716 116988
rect 65716 116932 65720 116988
rect 65656 116928 65720 116932
rect 65736 116988 65800 116992
rect 65736 116932 65740 116988
rect 65740 116932 65796 116988
rect 65796 116932 65800 116988
rect 65736 116928 65800 116932
rect 65816 116988 65880 116992
rect 65816 116932 65820 116988
rect 65820 116932 65876 116988
rect 65876 116932 65880 116988
rect 65816 116928 65880 116932
rect 65896 116988 65960 116992
rect 65896 116932 65900 116988
rect 65900 116932 65956 116988
rect 65956 116932 65960 116988
rect 65896 116928 65960 116932
rect 19576 116444 19640 116448
rect 19576 116388 19580 116444
rect 19580 116388 19636 116444
rect 19636 116388 19640 116444
rect 19576 116384 19640 116388
rect 19656 116444 19720 116448
rect 19656 116388 19660 116444
rect 19660 116388 19716 116444
rect 19716 116388 19720 116444
rect 19656 116384 19720 116388
rect 19736 116444 19800 116448
rect 19736 116388 19740 116444
rect 19740 116388 19796 116444
rect 19796 116388 19800 116444
rect 19736 116384 19800 116388
rect 19816 116444 19880 116448
rect 19816 116388 19820 116444
rect 19820 116388 19876 116444
rect 19876 116388 19880 116444
rect 19816 116384 19880 116388
rect 50296 116444 50360 116448
rect 50296 116388 50300 116444
rect 50300 116388 50356 116444
rect 50356 116388 50360 116444
rect 50296 116384 50360 116388
rect 50376 116444 50440 116448
rect 50376 116388 50380 116444
rect 50380 116388 50436 116444
rect 50436 116388 50440 116444
rect 50376 116384 50440 116388
rect 50456 116444 50520 116448
rect 50456 116388 50460 116444
rect 50460 116388 50516 116444
rect 50516 116388 50520 116444
rect 50456 116384 50520 116388
rect 50536 116444 50600 116448
rect 50536 116388 50540 116444
rect 50540 116388 50596 116444
rect 50596 116388 50600 116444
rect 50536 116384 50600 116388
rect 4216 115900 4280 115904
rect 4216 115844 4220 115900
rect 4220 115844 4276 115900
rect 4276 115844 4280 115900
rect 4216 115840 4280 115844
rect 4296 115900 4360 115904
rect 4296 115844 4300 115900
rect 4300 115844 4356 115900
rect 4356 115844 4360 115900
rect 4296 115840 4360 115844
rect 4376 115900 4440 115904
rect 4376 115844 4380 115900
rect 4380 115844 4436 115900
rect 4436 115844 4440 115900
rect 4376 115840 4440 115844
rect 4456 115900 4520 115904
rect 4456 115844 4460 115900
rect 4460 115844 4516 115900
rect 4516 115844 4520 115900
rect 4456 115840 4520 115844
rect 34936 115900 35000 115904
rect 34936 115844 34940 115900
rect 34940 115844 34996 115900
rect 34996 115844 35000 115900
rect 34936 115840 35000 115844
rect 35016 115900 35080 115904
rect 35016 115844 35020 115900
rect 35020 115844 35076 115900
rect 35076 115844 35080 115900
rect 35016 115840 35080 115844
rect 35096 115900 35160 115904
rect 35096 115844 35100 115900
rect 35100 115844 35156 115900
rect 35156 115844 35160 115900
rect 35096 115840 35160 115844
rect 35176 115900 35240 115904
rect 35176 115844 35180 115900
rect 35180 115844 35236 115900
rect 35236 115844 35240 115900
rect 35176 115840 35240 115844
rect 65656 115900 65720 115904
rect 65656 115844 65660 115900
rect 65660 115844 65716 115900
rect 65716 115844 65720 115900
rect 65656 115840 65720 115844
rect 65736 115900 65800 115904
rect 65736 115844 65740 115900
rect 65740 115844 65796 115900
rect 65796 115844 65800 115900
rect 65736 115840 65800 115844
rect 65816 115900 65880 115904
rect 65816 115844 65820 115900
rect 65820 115844 65876 115900
rect 65876 115844 65880 115900
rect 65816 115840 65880 115844
rect 65896 115900 65960 115904
rect 65896 115844 65900 115900
rect 65900 115844 65956 115900
rect 65956 115844 65960 115900
rect 65896 115840 65960 115844
rect 19576 115356 19640 115360
rect 19576 115300 19580 115356
rect 19580 115300 19636 115356
rect 19636 115300 19640 115356
rect 19576 115296 19640 115300
rect 19656 115356 19720 115360
rect 19656 115300 19660 115356
rect 19660 115300 19716 115356
rect 19716 115300 19720 115356
rect 19656 115296 19720 115300
rect 19736 115356 19800 115360
rect 19736 115300 19740 115356
rect 19740 115300 19796 115356
rect 19796 115300 19800 115356
rect 19736 115296 19800 115300
rect 19816 115356 19880 115360
rect 19816 115300 19820 115356
rect 19820 115300 19876 115356
rect 19876 115300 19880 115356
rect 19816 115296 19880 115300
rect 50296 115356 50360 115360
rect 50296 115300 50300 115356
rect 50300 115300 50356 115356
rect 50356 115300 50360 115356
rect 50296 115296 50360 115300
rect 50376 115356 50440 115360
rect 50376 115300 50380 115356
rect 50380 115300 50436 115356
rect 50436 115300 50440 115356
rect 50376 115296 50440 115300
rect 50456 115356 50520 115360
rect 50456 115300 50460 115356
rect 50460 115300 50516 115356
rect 50516 115300 50520 115356
rect 50456 115296 50520 115300
rect 50536 115356 50600 115360
rect 50536 115300 50540 115356
rect 50540 115300 50596 115356
rect 50596 115300 50600 115356
rect 50536 115296 50600 115300
rect 4216 114812 4280 114816
rect 4216 114756 4220 114812
rect 4220 114756 4276 114812
rect 4276 114756 4280 114812
rect 4216 114752 4280 114756
rect 4296 114812 4360 114816
rect 4296 114756 4300 114812
rect 4300 114756 4356 114812
rect 4356 114756 4360 114812
rect 4296 114752 4360 114756
rect 4376 114812 4440 114816
rect 4376 114756 4380 114812
rect 4380 114756 4436 114812
rect 4436 114756 4440 114812
rect 4376 114752 4440 114756
rect 4456 114812 4520 114816
rect 4456 114756 4460 114812
rect 4460 114756 4516 114812
rect 4516 114756 4520 114812
rect 4456 114752 4520 114756
rect 34936 114812 35000 114816
rect 34936 114756 34940 114812
rect 34940 114756 34996 114812
rect 34996 114756 35000 114812
rect 34936 114752 35000 114756
rect 35016 114812 35080 114816
rect 35016 114756 35020 114812
rect 35020 114756 35076 114812
rect 35076 114756 35080 114812
rect 35016 114752 35080 114756
rect 35096 114812 35160 114816
rect 35096 114756 35100 114812
rect 35100 114756 35156 114812
rect 35156 114756 35160 114812
rect 35096 114752 35160 114756
rect 35176 114812 35240 114816
rect 35176 114756 35180 114812
rect 35180 114756 35236 114812
rect 35236 114756 35240 114812
rect 35176 114752 35240 114756
rect 65656 114812 65720 114816
rect 65656 114756 65660 114812
rect 65660 114756 65716 114812
rect 65716 114756 65720 114812
rect 65656 114752 65720 114756
rect 65736 114812 65800 114816
rect 65736 114756 65740 114812
rect 65740 114756 65796 114812
rect 65796 114756 65800 114812
rect 65736 114752 65800 114756
rect 65816 114812 65880 114816
rect 65816 114756 65820 114812
rect 65820 114756 65876 114812
rect 65876 114756 65880 114812
rect 65816 114752 65880 114756
rect 65896 114812 65960 114816
rect 65896 114756 65900 114812
rect 65900 114756 65956 114812
rect 65956 114756 65960 114812
rect 65896 114752 65960 114756
rect 19576 114268 19640 114272
rect 19576 114212 19580 114268
rect 19580 114212 19636 114268
rect 19636 114212 19640 114268
rect 19576 114208 19640 114212
rect 19656 114268 19720 114272
rect 19656 114212 19660 114268
rect 19660 114212 19716 114268
rect 19716 114212 19720 114268
rect 19656 114208 19720 114212
rect 19736 114268 19800 114272
rect 19736 114212 19740 114268
rect 19740 114212 19796 114268
rect 19796 114212 19800 114268
rect 19736 114208 19800 114212
rect 19816 114268 19880 114272
rect 19816 114212 19820 114268
rect 19820 114212 19876 114268
rect 19876 114212 19880 114268
rect 19816 114208 19880 114212
rect 50296 114268 50360 114272
rect 50296 114212 50300 114268
rect 50300 114212 50356 114268
rect 50356 114212 50360 114268
rect 50296 114208 50360 114212
rect 50376 114268 50440 114272
rect 50376 114212 50380 114268
rect 50380 114212 50436 114268
rect 50436 114212 50440 114268
rect 50376 114208 50440 114212
rect 50456 114268 50520 114272
rect 50456 114212 50460 114268
rect 50460 114212 50516 114268
rect 50516 114212 50520 114268
rect 50456 114208 50520 114212
rect 50536 114268 50600 114272
rect 50536 114212 50540 114268
rect 50540 114212 50596 114268
rect 50596 114212 50600 114268
rect 50536 114208 50600 114212
rect 4216 113724 4280 113728
rect 4216 113668 4220 113724
rect 4220 113668 4276 113724
rect 4276 113668 4280 113724
rect 4216 113664 4280 113668
rect 4296 113724 4360 113728
rect 4296 113668 4300 113724
rect 4300 113668 4356 113724
rect 4356 113668 4360 113724
rect 4296 113664 4360 113668
rect 4376 113724 4440 113728
rect 4376 113668 4380 113724
rect 4380 113668 4436 113724
rect 4436 113668 4440 113724
rect 4376 113664 4440 113668
rect 4456 113724 4520 113728
rect 4456 113668 4460 113724
rect 4460 113668 4516 113724
rect 4516 113668 4520 113724
rect 4456 113664 4520 113668
rect 34936 113724 35000 113728
rect 34936 113668 34940 113724
rect 34940 113668 34996 113724
rect 34996 113668 35000 113724
rect 34936 113664 35000 113668
rect 35016 113724 35080 113728
rect 35016 113668 35020 113724
rect 35020 113668 35076 113724
rect 35076 113668 35080 113724
rect 35016 113664 35080 113668
rect 35096 113724 35160 113728
rect 35096 113668 35100 113724
rect 35100 113668 35156 113724
rect 35156 113668 35160 113724
rect 35096 113664 35160 113668
rect 35176 113724 35240 113728
rect 35176 113668 35180 113724
rect 35180 113668 35236 113724
rect 35236 113668 35240 113724
rect 35176 113664 35240 113668
rect 65656 113724 65720 113728
rect 65656 113668 65660 113724
rect 65660 113668 65716 113724
rect 65716 113668 65720 113724
rect 65656 113664 65720 113668
rect 65736 113724 65800 113728
rect 65736 113668 65740 113724
rect 65740 113668 65796 113724
rect 65796 113668 65800 113724
rect 65736 113664 65800 113668
rect 65816 113724 65880 113728
rect 65816 113668 65820 113724
rect 65820 113668 65876 113724
rect 65876 113668 65880 113724
rect 65816 113664 65880 113668
rect 65896 113724 65960 113728
rect 65896 113668 65900 113724
rect 65900 113668 65956 113724
rect 65956 113668 65960 113724
rect 65896 113664 65960 113668
rect 19576 113180 19640 113184
rect 19576 113124 19580 113180
rect 19580 113124 19636 113180
rect 19636 113124 19640 113180
rect 19576 113120 19640 113124
rect 19656 113180 19720 113184
rect 19656 113124 19660 113180
rect 19660 113124 19716 113180
rect 19716 113124 19720 113180
rect 19656 113120 19720 113124
rect 19736 113180 19800 113184
rect 19736 113124 19740 113180
rect 19740 113124 19796 113180
rect 19796 113124 19800 113180
rect 19736 113120 19800 113124
rect 19816 113180 19880 113184
rect 19816 113124 19820 113180
rect 19820 113124 19876 113180
rect 19876 113124 19880 113180
rect 19816 113120 19880 113124
rect 50296 113180 50360 113184
rect 50296 113124 50300 113180
rect 50300 113124 50356 113180
rect 50356 113124 50360 113180
rect 50296 113120 50360 113124
rect 50376 113180 50440 113184
rect 50376 113124 50380 113180
rect 50380 113124 50436 113180
rect 50436 113124 50440 113180
rect 50376 113120 50440 113124
rect 50456 113180 50520 113184
rect 50456 113124 50460 113180
rect 50460 113124 50516 113180
rect 50516 113124 50520 113180
rect 50456 113120 50520 113124
rect 50536 113180 50600 113184
rect 50536 113124 50540 113180
rect 50540 113124 50596 113180
rect 50596 113124 50600 113180
rect 50536 113120 50600 113124
rect 4216 112636 4280 112640
rect 4216 112580 4220 112636
rect 4220 112580 4276 112636
rect 4276 112580 4280 112636
rect 4216 112576 4280 112580
rect 4296 112636 4360 112640
rect 4296 112580 4300 112636
rect 4300 112580 4356 112636
rect 4356 112580 4360 112636
rect 4296 112576 4360 112580
rect 4376 112636 4440 112640
rect 4376 112580 4380 112636
rect 4380 112580 4436 112636
rect 4436 112580 4440 112636
rect 4376 112576 4440 112580
rect 4456 112636 4520 112640
rect 4456 112580 4460 112636
rect 4460 112580 4516 112636
rect 4516 112580 4520 112636
rect 4456 112576 4520 112580
rect 34936 112636 35000 112640
rect 34936 112580 34940 112636
rect 34940 112580 34996 112636
rect 34996 112580 35000 112636
rect 34936 112576 35000 112580
rect 35016 112636 35080 112640
rect 35016 112580 35020 112636
rect 35020 112580 35076 112636
rect 35076 112580 35080 112636
rect 35016 112576 35080 112580
rect 35096 112636 35160 112640
rect 35096 112580 35100 112636
rect 35100 112580 35156 112636
rect 35156 112580 35160 112636
rect 35096 112576 35160 112580
rect 35176 112636 35240 112640
rect 35176 112580 35180 112636
rect 35180 112580 35236 112636
rect 35236 112580 35240 112636
rect 35176 112576 35240 112580
rect 65656 112636 65720 112640
rect 65656 112580 65660 112636
rect 65660 112580 65716 112636
rect 65716 112580 65720 112636
rect 65656 112576 65720 112580
rect 65736 112636 65800 112640
rect 65736 112580 65740 112636
rect 65740 112580 65796 112636
rect 65796 112580 65800 112636
rect 65736 112576 65800 112580
rect 65816 112636 65880 112640
rect 65816 112580 65820 112636
rect 65820 112580 65876 112636
rect 65876 112580 65880 112636
rect 65816 112576 65880 112580
rect 65896 112636 65960 112640
rect 65896 112580 65900 112636
rect 65900 112580 65956 112636
rect 65956 112580 65960 112636
rect 65896 112576 65960 112580
rect 19576 112092 19640 112096
rect 19576 112036 19580 112092
rect 19580 112036 19636 112092
rect 19636 112036 19640 112092
rect 19576 112032 19640 112036
rect 19656 112092 19720 112096
rect 19656 112036 19660 112092
rect 19660 112036 19716 112092
rect 19716 112036 19720 112092
rect 19656 112032 19720 112036
rect 19736 112092 19800 112096
rect 19736 112036 19740 112092
rect 19740 112036 19796 112092
rect 19796 112036 19800 112092
rect 19736 112032 19800 112036
rect 19816 112092 19880 112096
rect 19816 112036 19820 112092
rect 19820 112036 19876 112092
rect 19876 112036 19880 112092
rect 19816 112032 19880 112036
rect 50296 112092 50360 112096
rect 50296 112036 50300 112092
rect 50300 112036 50356 112092
rect 50356 112036 50360 112092
rect 50296 112032 50360 112036
rect 50376 112092 50440 112096
rect 50376 112036 50380 112092
rect 50380 112036 50436 112092
rect 50436 112036 50440 112092
rect 50376 112032 50440 112036
rect 50456 112092 50520 112096
rect 50456 112036 50460 112092
rect 50460 112036 50516 112092
rect 50516 112036 50520 112092
rect 50456 112032 50520 112036
rect 50536 112092 50600 112096
rect 50536 112036 50540 112092
rect 50540 112036 50596 112092
rect 50596 112036 50600 112092
rect 50536 112032 50600 112036
rect 4216 111548 4280 111552
rect 4216 111492 4220 111548
rect 4220 111492 4276 111548
rect 4276 111492 4280 111548
rect 4216 111488 4280 111492
rect 4296 111548 4360 111552
rect 4296 111492 4300 111548
rect 4300 111492 4356 111548
rect 4356 111492 4360 111548
rect 4296 111488 4360 111492
rect 4376 111548 4440 111552
rect 4376 111492 4380 111548
rect 4380 111492 4436 111548
rect 4436 111492 4440 111548
rect 4376 111488 4440 111492
rect 4456 111548 4520 111552
rect 4456 111492 4460 111548
rect 4460 111492 4516 111548
rect 4516 111492 4520 111548
rect 4456 111488 4520 111492
rect 34936 111548 35000 111552
rect 34936 111492 34940 111548
rect 34940 111492 34996 111548
rect 34996 111492 35000 111548
rect 34936 111488 35000 111492
rect 35016 111548 35080 111552
rect 35016 111492 35020 111548
rect 35020 111492 35076 111548
rect 35076 111492 35080 111548
rect 35016 111488 35080 111492
rect 35096 111548 35160 111552
rect 35096 111492 35100 111548
rect 35100 111492 35156 111548
rect 35156 111492 35160 111548
rect 35096 111488 35160 111492
rect 35176 111548 35240 111552
rect 35176 111492 35180 111548
rect 35180 111492 35236 111548
rect 35236 111492 35240 111548
rect 35176 111488 35240 111492
rect 65656 111548 65720 111552
rect 65656 111492 65660 111548
rect 65660 111492 65716 111548
rect 65716 111492 65720 111548
rect 65656 111488 65720 111492
rect 65736 111548 65800 111552
rect 65736 111492 65740 111548
rect 65740 111492 65796 111548
rect 65796 111492 65800 111548
rect 65736 111488 65800 111492
rect 65816 111548 65880 111552
rect 65816 111492 65820 111548
rect 65820 111492 65876 111548
rect 65876 111492 65880 111548
rect 65816 111488 65880 111492
rect 65896 111548 65960 111552
rect 65896 111492 65900 111548
rect 65900 111492 65956 111548
rect 65956 111492 65960 111548
rect 65896 111488 65960 111492
rect 19576 111004 19640 111008
rect 19576 110948 19580 111004
rect 19580 110948 19636 111004
rect 19636 110948 19640 111004
rect 19576 110944 19640 110948
rect 19656 111004 19720 111008
rect 19656 110948 19660 111004
rect 19660 110948 19716 111004
rect 19716 110948 19720 111004
rect 19656 110944 19720 110948
rect 19736 111004 19800 111008
rect 19736 110948 19740 111004
rect 19740 110948 19796 111004
rect 19796 110948 19800 111004
rect 19736 110944 19800 110948
rect 19816 111004 19880 111008
rect 19816 110948 19820 111004
rect 19820 110948 19876 111004
rect 19876 110948 19880 111004
rect 19816 110944 19880 110948
rect 50296 111004 50360 111008
rect 50296 110948 50300 111004
rect 50300 110948 50356 111004
rect 50356 110948 50360 111004
rect 50296 110944 50360 110948
rect 50376 111004 50440 111008
rect 50376 110948 50380 111004
rect 50380 110948 50436 111004
rect 50436 110948 50440 111004
rect 50376 110944 50440 110948
rect 50456 111004 50520 111008
rect 50456 110948 50460 111004
rect 50460 110948 50516 111004
rect 50516 110948 50520 111004
rect 50456 110944 50520 110948
rect 50536 111004 50600 111008
rect 50536 110948 50540 111004
rect 50540 110948 50596 111004
rect 50596 110948 50600 111004
rect 50536 110944 50600 110948
rect 4216 110460 4280 110464
rect 4216 110404 4220 110460
rect 4220 110404 4276 110460
rect 4276 110404 4280 110460
rect 4216 110400 4280 110404
rect 4296 110460 4360 110464
rect 4296 110404 4300 110460
rect 4300 110404 4356 110460
rect 4356 110404 4360 110460
rect 4296 110400 4360 110404
rect 4376 110460 4440 110464
rect 4376 110404 4380 110460
rect 4380 110404 4436 110460
rect 4436 110404 4440 110460
rect 4376 110400 4440 110404
rect 4456 110460 4520 110464
rect 4456 110404 4460 110460
rect 4460 110404 4516 110460
rect 4516 110404 4520 110460
rect 4456 110400 4520 110404
rect 34936 110460 35000 110464
rect 34936 110404 34940 110460
rect 34940 110404 34996 110460
rect 34996 110404 35000 110460
rect 34936 110400 35000 110404
rect 35016 110460 35080 110464
rect 35016 110404 35020 110460
rect 35020 110404 35076 110460
rect 35076 110404 35080 110460
rect 35016 110400 35080 110404
rect 35096 110460 35160 110464
rect 35096 110404 35100 110460
rect 35100 110404 35156 110460
rect 35156 110404 35160 110460
rect 35096 110400 35160 110404
rect 35176 110460 35240 110464
rect 35176 110404 35180 110460
rect 35180 110404 35236 110460
rect 35236 110404 35240 110460
rect 35176 110400 35240 110404
rect 65656 110460 65720 110464
rect 65656 110404 65660 110460
rect 65660 110404 65716 110460
rect 65716 110404 65720 110460
rect 65656 110400 65720 110404
rect 65736 110460 65800 110464
rect 65736 110404 65740 110460
rect 65740 110404 65796 110460
rect 65796 110404 65800 110460
rect 65736 110400 65800 110404
rect 65816 110460 65880 110464
rect 65816 110404 65820 110460
rect 65820 110404 65876 110460
rect 65876 110404 65880 110460
rect 65816 110400 65880 110404
rect 65896 110460 65960 110464
rect 65896 110404 65900 110460
rect 65900 110404 65956 110460
rect 65956 110404 65960 110460
rect 65896 110400 65960 110404
rect 19576 109916 19640 109920
rect 19576 109860 19580 109916
rect 19580 109860 19636 109916
rect 19636 109860 19640 109916
rect 19576 109856 19640 109860
rect 19656 109916 19720 109920
rect 19656 109860 19660 109916
rect 19660 109860 19716 109916
rect 19716 109860 19720 109916
rect 19656 109856 19720 109860
rect 19736 109916 19800 109920
rect 19736 109860 19740 109916
rect 19740 109860 19796 109916
rect 19796 109860 19800 109916
rect 19736 109856 19800 109860
rect 19816 109916 19880 109920
rect 19816 109860 19820 109916
rect 19820 109860 19876 109916
rect 19876 109860 19880 109916
rect 19816 109856 19880 109860
rect 50296 109916 50360 109920
rect 50296 109860 50300 109916
rect 50300 109860 50356 109916
rect 50356 109860 50360 109916
rect 50296 109856 50360 109860
rect 50376 109916 50440 109920
rect 50376 109860 50380 109916
rect 50380 109860 50436 109916
rect 50436 109860 50440 109916
rect 50376 109856 50440 109860
rect 50456 109916 50520 109920
rect 50456 109860 50460 109916
rect 50460 109860 50516 109916
rect 50516 109860 50520 109916
rect 50456 109856 50520 109860
rect 50536 109916 50600 109920
rect 50536 109860 50540 109916
rect 50540 109860 50596 109916
rect 50596 109860 50600 109916
rect 50536 109856 50600 109860
rect 4216 109372 4280 109376
rect 4216 109316 4220 109372
rect 4220 109316 4276 109372
rect 4276 109316 4280 109372
rect 4216 109312 4280 109316
rect 4296 109372 4360 109376
rect 4296 109316 4300 109372
rect 4300 109316 4356 109372
rect 4356 109316 4360 109372
rect 4296 109312 4360 109316
rect 4376 109372 4440 109376
rect 4376 109316 4380 109372
rect 4380 109316 4436 109372
rect 4436 109316 4440 109372
rect 4376 109312 4440 109316
rect 4456 109372 4520 109376
rect 4456 109316 4460 109372
rect 4460 109316 4516 109372
rect 4516 109316 4520 109372
rect 4456 109312 4520 109316
rect 34936 109372 35000 109376
rect 34936 109316 34940 109372
rect 34940 109316 34996 109372
rect 34996 109316 35000 109372
rect 34936 109312 35000 109316
rect 35016 109372 35080 109376
rect 35016 109316 35020 109372
rect 35020 109316 35076 109372
rect 35076 109316 35080 109372
rect 35016 109312 35080 109316
rect 35096 109372 35160 109376
rect 35096 109316 35100 109372
rect 35100 109316 35156 109372
rect 35156 109316 35160 109372
rect 35096 109312 35160 109316
rect 35176 109372 35240 109376
rect 35176 109316 35180 109372
rect 35180 109316 35236 109372
rect 35236 109316 35240 109372
rect 35176 109312 35240 109316
rect 65656 109372 65720 109376
rect 65656 109316 65660 109372
rect 65660 109316 65716 109372
rect 65716 109316 65720 109372
rect 65656 109312 65720 109316
rect 65736 109372 65800 109376
rect 65736 109316 65740 109372
rect 65740 109316 65796 109372
rect 65796 109316 65800 109372
rect 65736 109312 65800 109316
rect 65816 109372 65880 109376
rect 65816 109316 65820 109372
rect 65820 109316 65876 109372
rect 65876 109316 65880 109372
rect 65816 109312 65880 109316
rect 65896 109372 65960 109376
rect 65896 109316 65900 109372
rect 65900 109316 65956 109372
rect 65956 109316 65960 109372
rect 65896 109312 65960 109316
rect 19576 108828 19640 108832
rect 19576 108772 19580 108828
rect 19580 108772 19636 108828
rect 19636 108772 19640 108828
rect 19576 108768 19640 108772
rect 19656 108828 19720 108832
rect 19656 108772 19660 108828
rect 19660 108772 19716 108828
rect 19716 108772 19720 108828
rect 19656 108768 19720 108772
rect 19736 108828 19800 108832
rect 19736 108772 19740 108828
rect 19740 108772 19796 108828
rect 19796 108772 19800 108828
rect 19736 108768 19800 108772
rect 19816 108828 19880 108832
rect 19816 108772 19820 108828
rect 19820 108772 19876 108828
rect 19876 108772 19880 108828
rect 19816 108768 19880 108772
rect 50296 108828 50360 108832
rect 50296 108772 50300 108828
rect 50300 108772 50356 108828
rect 50356 108772 50360 108828
rect 50296 108768 50360 108772
rect 50376 108828 50440 108832
rect 50376 108772 50380 108828
rect 50380 108772 50436 108828
rect 50436 108772 50440 108828
rect 50376 108768 50440 108772
rect 50456 108828 50520 108832
rect 50456 108772 50460 108828
rect 50460 108772 50516 108828
rect 50516 108772 50520 108828
rect 50456 108768 50520 108772
rect 50536 108828 50600 108832
rect 50536 108772 50540 108828
rect 50540 108772 50596 108828
rect 50596 108772 50600 108828
rect 50536 108768 50600 108772
rect 4216 108284 4280 108288
rect 4216 108228 4220 108284
rect 4220 108228 4276 108284
rect 4276 108228 4280 108284
rect 4216 108224 4280 108228
rect 4296 108284 4360 108288
rect 4296 108228 4300 108284
rect 4300 108228 4356 108284
rect 4356 108228 4360 108284
rect 4296 108224 4360 108228
rect 4376 108284 4440 108288
rect 4376 108228 4380 108284
rect 4380 108228 4436 108284
rect 4436 108228 4440 108284
rect 4376 108224 4440 108228
rect 4456 108284 4520 108288
rect 4456 108228 4460 108284
rect 4460 108228 4516 108284
rect 4516 108228 4520 108284
rect 4456 108224 4520 108228
rect 34936 108284 35000 108288
rect 34936 108228 34940 108284
rect 34940 108228 34996 108284
rect 34996 108228 35000 108284
rect 34936 108224 35000 108228
rect 35016 108284 35080 108288
rect 35016 108228 35020 108284
rect 35020 108228 35076 108284
rect 35076 108228 35080 108284
rect 35016 108224 35080 108228
rect 35096 108284 35160 108288
rect 35096 108228 35100 108284
rect 35100 108228 35156 108284
rect 35156 108228 35160 108284
rect 35096 108224 35160 108228
rect 35176 108284 35240 108288
rect 35176 108228 35180 108284
rect 35180 108228 35236 108284
rect 35236 108228 35240 108284
rect 35176 108224 35240 108228
rect 65656 108284 65720 108288
rect 65656 108228 65660 108284
rect 65660 108228 65716 108284
rect 65716 108228 65720 108284
rect 65656 108224 65720 108228
rect 65736 108284 65800 108288
rect 65736 108228 65740 108284
rect 65740 108228 65796 108284
rect 65796 108228 65800 108284
rect 65736 108224 65800 108228
rect 65816 108284 65880 108288
rect 65816 108228 65820 108284
rect 65820 108228 65876 108284
rect 65876 108228 65880 108284
rect 65816 108224 65880 108228
rect 65896 108284 65960 108288
rect 65896 108228 65900 108284
rect 65900 108228 65956 108284
rect 65956 108228 65960 108284
rect 65896 108224 65960 108228
rect 19576 107740 19640 107744
rect 19576 107684 19580 107740
rect 19580 107684 19636 107740
rect 19636 107684 19640 107740
rect 19576 107680 19640 107684
rect 19656 107740 19720 107744
rect 19656 107684 19660 107740
rect 19660 107684 19716 107740
rect 19716 107684 19720 107740
rect 19656 107680 19720 107684
rect 19736 107740 19800 107744
rect 19736 107684 19740 107740
rect 19740 107684 19796 107740
rect 19796 107684 19800 107740
rect 19736 107680 19800 107684
rect 19816 107740 19880 107744
rect 19816 107684 19820 107740
rect 19820 107684 19876 107740
rect 19876 107684 19880 107740
rect 19816 107680 19880 107684
rect 50296 107740 50360 107744
rect 50296 107684 50300 107740
rect 50300 107684 50356 107740
rect 50356 107684 50360 107740
rect 50296 107680 50360 107684
rect 50376 107740 50440 107744
rect 50376 107684 50380 107740
rect 50380 107684 50436 107740
rect 50436 107684 50440 107740
rect 50376 107680 50440 107684
rect 50456 107740 50520 107744
rect 50456 107684 50460 107740
rect 50460 107684 50516 107740
rect 50516 107684 50520 107740
rect 50456 107680 50520 107684
rect 50536 107740 50600 107744
rect 50536 107684 50540 107740
rect 50540 107684 50596 107740
rect 50596 107684 50600 107740
rect 50536 107680 50600 107684
rect 4216 107196 4280 107200
rect 4216 107140 4220 107196
rect 4220 107140 4276 107196
rect 4276 107140 4280 107196
rect 4216 107136 4280 107140
rect 4296 107196 4360 107200
rect 4296 107140 4300 107196
rect 4300 107140 4356 107196
rect 4356 107140 4360 107196
rect 4296 107136 4360 107140
rect 4376 107196 4440 107200
rect 4376 107140 4380 107196
rect 4380 107140 4436 107196
rect 4436 107140 4440 107196
rect 4376 107136 4440 107140
rect 4456 107196 4520 107200
rect 4456 107140 4460 107196
rect 4460 107140 4516 107196
rect 4516 107140 4520 107196
rect 4456 107136 4520 107140
rect 34936 107196 35000 107200
rect 34936 107140 34940 107196
rect 34940 107140 34996 107196
rect 34996 107140 35000 107196
rect 34936 107136 35000 107140
rect 35016 107196 35080 107200
rect 35016 107140 35020 107196
rect 35020 107140 35076 107196
rect 35076 107140 35080 107196
rect 35016 107136 35080 107140
rect 35096 107196 35160 107200
rect 35096 107140 35100 107196
rect 35100 107140 35156 107196
rect 35156 107140 35160 107196
rect 35096 107136 35160 107140
rect 35176 107196 35240 107200
rect 35176 107140 35180 107196
rect 35180 107140 35236 107196
rect 35236 107140 35240 107196
rect 35176 107136 35240 107140
rect 65656 107196 65720 107200
rect 65656 107140 65660 107196
rect 65660 107140 65716 107196
rect 65716 107140 65720 107196
rect 65656 107136 65720 107140
rect 65736 107196 65800 107200
rect 65736 107140 65740 107196
rect 65740 107140 65796 107196
rect 65796 107140 65800 107196
rect 65736 107136 65800 107140
rect 65816 107196 65880 107200
rect 65816 107140 65820 107196
rect 65820 107140 65876 107196
rect 65876 107140 65880 107196
rect 65816 107136 65880 107140
rect 65896 107196 65960 107200
rect 65896 107140 65900 107196
rect 65900 107140 65956 107196
rect 65956 107140 65960 107196
rect 65896 107136 65960 107140
rect 19576 106652 19640 106656
rect 19576 106596 19580 106652
rect 19580 106596 19636 106652
rect 19636 106596 19640 106652
rect 19576 106592 19640 106596
rect 19656 106652 19720 106656
rect 19656 106596 19660 106652
rect 19660 106596 19716 106652
rect 19716 106596 19720 106652
rect 19656 106592 19720 106596
rect 19736 106652 19800 106656
rect 19736 106596 19740 106652
rect 19740 106596 19796 106652
rect 19796 106596 19800 106652
rect 19736 106592 19800 106596
rect 19816 106652 19880 106656
rect 19816 106596 19820 106652
rect 19820 106596 19876 106652
rect 19876 106596 19880 106652
rect 19816 106592 19880 106596
rect 50296 106652 50360 106656
rect 50296 106596 50300 106652
rect 50300 106596 50356 106652
rect 50356 106596 50360 106652
rect 50296 106592 50360 106596
rect 50376 106652 50440 106656
rect 50376 106596 50380 106652
rect 50380 106596 50436 106652
rect 50436 106596 50440 106652
rect 50376 106592 50440 106596
rect 50456 106652 50520 106656
rect 50456 106596 50460 106652
rect 50460 106596 50516 106652
rect 50516 106596 50520 106652
rect 50456 106592 50520 106596
rect 50536 106652 50600 106656
rect 50536 106596 50540 106652
rect 50540 106596 50596 106652
rect 50596 106596 50600 106652
rect 50536 106592 50600 106596
rect 4216 106108 4280 106112
rect 4216 106052 4220 106108
rect 4220 106052 4276 106108
rect 4276 106052 4280 106108
rect 4216 106048 4280 106052
rect 4296 106108 4360 106112
rect 4296 106052 4300 106108
rect 4300 106052 4356 106108
rect 4356 106052 4360 106108
rect 4296 106048 4360 106052
rect 4376 106108 4440 106112
rect 4376 106052 4380 106108
rect 4380 106052 4436 106108
rect 4436 106052 4440 106108
rect 4376 106048 4440 106052
rect 4456 106108 4520 106112
rect 4456 106052 4460 106108
rect 4460 106052 4516 106108
rect 4516 106052 4520 106108
rect 4456 106048 4520 106052
rect 34936 106108 35000 106112
rect 34936 106052 34940 106108
rect 34940 106052 34996 106108
rect 34996 106052 35000 106108
rect 34936 106048 35000 106052
rect 35016 106108 35080 106112
rect 35016 106052 35020 106108
rect 35020 106052 35076 106108
rect 35076 106052 35080 106108
rect 35016 106048 35080 106052
rect 35096 106108 35160 106112
rect 35096 106052 35100 106108
rect 35100 106052 35156 106108
rect 35156 106052 35160 106108
rect 35096 106048 35160 106052
rect 35176 106108 35240 106112
rect 35176 106052 35180 106108
rect 35180 106052 35236 106108
rect 35236 106052 35240 106108
rect 35176 106048 35240 106052
rect 65656 106108 65720 106112
rect 65656 106052 65660 106108
rect 65660 106052 65716 106108
rect 65716 106052 65720 106108
rect 65656 106048 65720 106052
rect 65736 106108 65800 106112
rect 65736 106052 65740 106108
rect 65740 106052 65796 106108
rect 65796 106052 65800 106108
rect 65736 106048 65800 106052
rect 65816 106108 65880 106112
rect 65816 106052 65820 106108
rect 65820 106052 65876 106108
rect 65876 106052 65880 106108
rect 65816 106048 65880 106052
rect 65896 106108 65960 106112
rect 65896 106052 65900 106108
rect 65900 106052 65956 106108
rect 65956 106052 65960 106108
rect 65896 106048 65960 106052
rect 19576 105564 19640 105568
rect 19576 105508 19580 105564
rect 19580 105508 19636 105564
rect 19636 105508 19640 105564
rect 19576 105504 19640 105508
rect 19656 105564 19720 105568
rect 19656 105508 19660 105564
rect 19660 105508 19716 105564
rect 19716 105508 19720 105564
rect 19656 105504 19720 105508
rect 19736 105564 19800 105568
rect 19736 105508 19740 105564
rect 19740 105508 19796 105564
rect 19796 105508 19800 105564
rect 19736 105504 19800 105508
rect 19816 105564 19880 105568
rect 19816 105508 19820 105564
rect 19820 105508 19876 105564
rect 19876 105508 19880 105564
rect 19816 105504 19880 105508
rect 50296 105564 50360 105568
rect 50296 105508 50300 105564
rect 50300 105508 50356 105564
rect 50356 105508 50360 105564
rect 50296 105504 50360 105508
rect 50376 105564 50440 105568
rect 50376 105508 50380 105564
rect 50380 105508 50436 105564
rect 50436 105508 50440 105564
rect 50376 105504 50440 105508
rect 50456 105564 50520 105568
rect 50456 105508 50460 105564
rect 50460 105508 50516 105564
rect 50516 105508 50520 105564
rect 50456 105504 50520 105508
rect 50536 105564 50600 105568
rect 50536 105508 50540 105564
rect 50540 105508 50596 105564
rect 50596 105508 50600 105564
rect 50536 105504 50600 105508
rect 4216 105020 4280 105024
rect 4216 104964 4220 105020
rect 4220 104964 4276 105020
rect 4276 104964 4280 105020
rect 4216 104960 4280 104964
rect 4296 105020 4360 105024
rect 4296 104964 4300 105020
rect 4300 104964 4356 105020
rect 4356 104964 4360 105020
rect 4296 104960 4360 104964
rect 4376 105020 4440 105024
rect 4376 104964 4380 105020
rect 4380 104964 4436 105020
rect 4436 104964 4440 105020
rect 4376 104960 4440 104964
rect 4456 105020 4520 105024
rect 4456 104964 4460 105020
rect 4460 104964 4516 105020
rect 4516 104964 4520 105020
rect 4456 104960 4520 104964
rect 34936 105020 35000 105024
rect 34936 104964 34940 105020
rect 34940 104964 34996 105020
rect 34996 104964 35000 105020
rect 34936 104960 35000 104964
rect 35016 105020 35080 105024
rect 35016 104964 35020 105020
rect 35020 104964 35076 105020
rect 35076 104964 35080 105020
rect 35016 104960 35080 104964
rect 35096 105020 35160 105024
rect 35096 104964 35100 105020
rect 35100 104964 35156 105020
rect 35156 104964 35160 105020
rect 35096 104960 35160 104964
rect 35176 105020 35240 105024
rect 35176 104964 35180 105020
rect 35180 104964 35236 105020
rect 35236 104964 35240 105020
rect 35176 104960 35240 104964
rect 65656 105020 65720 105024
rect 65656 104964 65660 105020
rect 65660 104964 65716 105020
rect 65716 104964 65720 105020
rect 65656 104960 65720 104964
rect 65736 105020 65800 105024
rect 65736 104964 65740 105020
rect 65740 104964 65796 105020
rect 65796 104964 65800 105020
rect 65736 104960 65800 104964
rect 65816 105020 65880 105024
rect 65816 104964 65820 105020
rect 65820 104964 65876 105020
rect 65876 104964 65880 105020
rect 65816 104960 65880 104964
rect 65896 105020 65960 105024
rect 65896 104964 65900 105020
rect 65900 104964 65956 105020
rect 65956 104964 65960 105020
rect 65896 104960 65960 104964
rect 19576 104476 19640 104480
rect 19576 104420 19580 104476
rect 19580 104420 19636 104476
rect 19636 104420 19640 104476
rect 19576 104416 19640 104420
rect 19656 104476 19720 104480
rect 19656 104420 19660 104476
rect 19660 104420 19716 104476
rect 19716 104420 19720 104476
rect 19656 104416 19720 104420
rect 19736 104476 19800 104480
rect 19736 104420 19740 104476
rect 19740 104420 19796 104476
rect 19796 104420 19800 104476
rect 19736 104416 19800 104420
rect 19816 104476 19880 104480
rect 19816 104420 19820 104476
rect 19820 104420 19876 104476
rect 19876 104420 19880 104476
rect 19816 104416 19880 104420
rect 50296 104476 50360 104480
rect 50296 104420 50300 104476
rect 50300 104420 50356 104476
rect 50356 104420 50360 104476
rect 50296 104416 50360 104420
rect 50376 104476 50440 104480
rect 50376 104420 50380 104476
rect 50380 104420 50436 104476
rect 50436 104420 50440 104476
rect 50376 104416 50440 104420
rect 50456 104476 50520 104480
rect 50456 104420 50460 104476
rect 50460 104420 50516 104476
rect 50516 104420 50520 104476
rect 50456 104416 50520 104420
rect 50536 104476 50600 104480
rect 50536 104420 50540 104476
rect 50540 104420 50596 104476
rect 50596 104420 50600 104476
rect 50536 104416 50600 104420
rect 4216 103932 4280 103936
rect 4216 103876 4220 103932
rect 4220 103876 4276 103932
rect 4276 103876 4280 103932
rect 4216 103872 4280 103876
rect 4296 103932 4360 103936
rect 4296 103876 4300 103932
rect 4300 103876 4356 103932
rect 4356 103876 4360 103932
rect 4296 103872 4360 103876
rect 4376 103932 4440 103936
rect 4376 103876 4380 103932
rect 4380 103876 4436 103932
rect 4436 103876 4440 103932
rect 4376 103872 4440 103876
rect 4456 103932 4520 103936
rect 4456 103876 4460 103932
rect 4460 103876 4516 103932
rect 4516 103876 4520 103932
rect 4456 103872 4520 103876
rect 34936 103932 35000 103936
rect 34936 103876 34940 103932
rect 34940 103876 34996 103932
rect 34996 103876 35000 103932
rect 34936 103872 35000 103876
rect 35016 103932 35080 103936
rect 35016 103876 35020 103932
rect 35020 103876 35076 103932
rect 35076 103876 35080 103932
rect 35016 103872 35080 103876
rect 35096 103932 35160 103936
rect 35096 103876 35100 103932
rect 35100 103876 35156 103932
rect 35156 103876 35160 103932
rect 35096 103872 35160 103876
rect 35176 103932 35240 103936
rect 35176 103876 35180 103932
rect 35180 103876 35236 103932
rect 35236 103876 35240 103932
rect 35176 103872 35240 103876
rect 65656 103932 65720 103936
rect 65656 103876 65660 103932
rect 65660 103876 65716 103932
rect 65716 103876 65720 103932
rect 65656 103872 65720 103876
rect 65736 103932 65800 103936
rect 65736 103876 65740 103932
rect 65740 103876 65796 103932
rect 65796 103876 65800 103932
rect 65736 103872 65800 103876
rect 65816 103932 65880 103936
rect 65816 103876 65820 103932
rect 65820 103876 65876 103932
rect 65876 103876 65880 103932
rect 65816 103872 65880 103876
rect 65896 103932 65960 103936
rect 65896 103876 65900 103932
rect 65900 103876 65956 103932
rect 65956 103876 65960 103932
rect 65896 103872 65960 103876
rect 19576 103388 19640 103392
rect 19576 103332 19580 103388
rect 19580 103332 19636 103388
rect 19636 103332 19640 103388
rect 19576 103328 19640 103332
rect 19656 103388 19720 103392
rect 19656 103332 19660 103388
rect 19660 103332 19716 103388
rect 19716 103332 19720 103388
rect 19656 103328 19720 103332
rect 19736 103388 19800 103392
rect 19736 103332 19740 103388
rect 19740 103332 19796 103388
rect 19796 103332 19800 103388
rect 19736 103328 19800 103332
rect 19816 103388 19880 103392
rect 19816 103332 19820 103388
rect 19820 103332 19876 103388
rect 19876 103332 19880 103388
rect 19816 103328 19880 103332
rect 50296 103388 50360 103392
rect 50296 103332 50300 103388
rect 50300 103332 50356 103388
rect 50356 103332 50360 103388
rect 50296 103328 50360 103332
rect 50376 103388 50440 103392
rect 50376 103332 50380 103388
rect 50380 103332 50436 103388
rect 50436 103332 50440 103388
rect 50376 103328 50440 103332
rect 50456 103388 50520 103392
rect 50456 103332 50460 103388
rect 50460 103332 50516 103388
rect 50516 103332 50520 103388
rect 50456 103328 50520 103332
rect 50536 103388 50600 103392
rect 50536 103332 50540 103388
rect 50540 103332 50596 103388
rect 50596 103332 50600 103388
rect 50536 103328 50600 103332
rect 4216 102844 4280 102848
rect 4216 102788 4220 102844
rect 4220 102788 4276 102844
rect 4276 102788 4280 102844
rect 4216 102784 4280 102788
rect 4296 102844 4360 102848
rect 4296 102788 4300 102844
rect 4300 102788 4356 102844
rect 4356 102788 4360 102844
rect 4296 102784 4360 102788
rect 4376 102844 4440 102848
rect 4376 102788 4380 102844
rect 4380 102788 4436 102844
rect 4436 102788 4440 102844
rect 4376 102784 4440 102788
rect 4456 102844 4520 102848
rect 4456 102788 4460 102844
rect 4460 102788 4516 102844
rect 4516 102788 4520 102844
rect 4456 102784 4520 102788
rect 34936 102844 35000 102848
rect 34936 102788 34940 102844
rect 34940 102788 34996 102844
rect 34996 102788 35000 102844
rect 34936 102784 35000 102788
rect 35016 102844 35080 102848
rect 35016 102788 35020 102844
rect 35020 102788 35076 102844
rect 35076 102788 35080 102844
rect 35016 102784 35080 102788
rect 35096 102844 35160 102848
rect 35096 102788 35100 102844
rect 35100 102788 35156 102844
rect 35156 102788 35160 102844
rect 35096 102784 35160 102788
rect 35176 102844 35240 102848
rect 35176 102788 35180 102844
rect 35180 102788 35236 102844
rect 35236 102788 35240 102844
rect 35176 102784 35240 102788
rect 65656 102844 65720 102848
rect 65656 102788 65660 102844
rect 65660 102788 65716 102844
rect 65716 102788 65720 102844
rect 65656 102784 65720 102788
rect 65736 102844 65800 102848
rect 65736 102788 65740 102844
rect 65740 102788 65796 102844
rect 65796 102788 65800 102844
rect 65736 102784 65800 102788
rect 65816 102844 65880 102848
rect 65816 102788 65820 102844
rect 65820 102788 65876 102844
rect 65876 102788 65880 102844
rect 65816 102784 65880 102788
rect 65896 102844 65960 102848
rect 65896 102788 65900 102844
rect 65900 102788 65956 102844
rect 65956 102788 65960 102844
rect 65896 102784 65960 102788
rect 19576 102300 19640 102304
rect 19576 102244 19580 102300
rect 19580 102244 19636 102300
rect 19636 102244 19640 102300
rect 19576 102240 19640 102244
rect 19656 102300 19720 102304
rect 19656 102244 19660 102300
rect 19660 102244 19716 102300
rect 19716 102244 19720 102300
rect 19656 102240 19720 102244
rect 19736 102300 19800 102304
rect 19736 102244 19740 102300
rect 19740 102244 19796 102300
rect 19796 102244 19800 102300
rect 19736 102240 19800 102244
rect 19816 102300 19880 102304
rect 19816 102244 19820 102300
rect 19820 102244 19876 102300
rect 19876 102244 19880 102300
rect 19816 102240 19880 102244
rect 50296 102300 50360 102304
rect 50296 102244 50300 102300
rect 50300 102244 50356 102300
rect 50356 102244 50360 102300
rect 50296 102240 50360 102244
rect 50376 102300 50440 102304
rect 50376 102244 50380 102300
rect 50380 102244 50436 102300
rect 50436 102244 50440 102300
rect 50376 102240 50440 102244
rect 50456 102300 50520 102304
rect 50456 102244 50460 102300
rect 50460 102244 50516 102300
rect 50516 102244 50520 102300
rect 50456 102240 50520 102244
rect 50536 102300 50600 102304
rect 50536 102244 50540 102300
rect 50540 102244 50596 102300
rect 50596 102244 50600 102300
rect 50536 102240 50600 102244
rect 4216 101756 4280 101760
rect 4216 101700 4220 101756
rect 4220 101700 4276 101756
rect 4276 101700 4280 101756
rect 4216 101696 4280 101700
rect 4296 101756 4360 101760
rect 4296 101700 4300 101756
rect 4300 101700 4356 101756
rect 4356 101700 4360 101756
rect 4296 101696 4360 101700
rect 4376 101756 4440 101760
rect 4376 101700 4380 101756
rect 4380 101700 4436 101756
rect 4436 101700 4440 101756
rect 4376 101696 4440 101700
rect 4456 101756 4520 101760
rect 4456 101700 4460 101756
rect 4460 101700 4516 101756
rect 4516 101700 4520 101756
rect 4456 101696 4520 101700
rect 34936 101756 35000 101760
rect 34936 101700 34940 101756
rect 34940 101700 34996 101756
rect 34996 101700 35000 101756
rect 34936 101696 35000 101700
rect 35016 101756 35080 101760
rect 35016 101700 35020 101756
rect 35020 101700 35076 101756
rect 35076 101700 35080 101756
rect 35016 101696 35080 101700
rect 35096 101756 35160 101760
rect 35096 101700 35100 101756
rect 35100 101700 35156 101756
rect 35156 101700 35160 101756
rect 35096 101696 35160 101700
rect 35176 101756 35240 101760
rect 35176 101700 35180 101756
rect 35180 101700 35236 101756
rect 35236 101700 35240 101756
rect 35176 101696 35240 101700
rect 65656 101756 65720 101760
rect 65656 101700 65660 101756
rect 65660 101700 65716 101756
rect 65716 101700 65720 101756
rect 65656 101696 65720 101700
rect 65736 101756 65800 101760
rect 65736 101700 65740 101756
rect 65740 101700 65796 101756
rect 65796 101700 65800 101756
rect 65736 101696 65800 101700
rect 65816 101756 65880 101760
rect 65816 101700 65820 101756
rect 65820 101700 65876 101756
rect 65876 101700 65880 101756
rect 65816 101696 65880 101700
rect 65896 101756 65960 101760
rect 65896 101700 65900 101756
rect 65900 101700 65956 101756
rect 65956 101700 65960 101756
rect 65896 101696 65960 101700
rect 19576 101212 19640 101216
rect 19576 101156 19580 101212
rect 19580 101156 19636 101212
rect 19636 101156 19640 101212
rect 19576 101152 19640 101156
rect 19656 101212 19720 101216
rect 19656 101156 19660 101212
rect 19660 101156 19716 101212
rect 19716 101156 19720 101212
rect 19656 101152 19720 101156
rect 19736 101212 19800 101216
rect 19736 101156 19740 101212
rect 19740 101156 19796 101212
rect 19796 101156 19800 101212
rect 19736 101152 19800 101156
rect 19816 101212 19880 101216
rect 19816 101156 19820 101212
rect 19820 101156 19876 101212
rect 19876 101156 19880 101212
rect 19816 101152 19880 101156
rect 50296 101212 50360 101216
rect 50296 101156 50300 101212
rect 50300 101156 50356 101212
rect 50356 101156 50360 101212
rect 50296 101152 50360 101156
rect 50376 101212 50440 101216
rect 50376 101156 50380 101212
rect 50380 101156 50436 101212
rect 50436 101156 50440 101212
rect 50376 101152 50440 101156
rect 50456 101212 50520 101216
rect 50456 101156 50460 101212
rect 50460 101156 50516 101212
rect 50516 101156 50520 101212
rect 50456 101152 50520 101156
rect 50536 101212 50600 101216
rect 50536 101156 50540 101212
rect 50540 101156 50596 101212
rect 50596 101156 50600 101212
rect 50536 101152 50600 101156
rect 4216 100668 4280 100672
rect 4216 100612 4220 100668
rect 4220 100612 4276 100668
rect 4276 100612 4280 100668
rect 4216 100608 4280 100612
rect 4296 100668 4360 100672
rect 4296 100612 4300 100668
rect 4300 100612 4356 100668
rect 4356 100612 4360 100668
rect 4296 100608 4360 100612
rect 4376 100668 4440 100672
rect 4376 100612 4380 100668
rect 4380 100612 4436 100668
rect 4436 100612 4440 100668
rect 4376 100608 4440 100612
rect 4456 100668 4520 100672
rect 4456 100612 4460 100668
rect 4460 100612 4516 100668
rect 4516 100612 4520 100668
rect 4456 100608 4520 100612
rect 34936 100668 35000 100672
rect 34936 100612 34940 100668
rect 34940 100612 34996 100668
rect 34996 100612 35000 100668
rect 34936 100608 35000 100612
rect 35016 100668 35080 100672
rect 35016 100612 35020 100668
rect 35020 100612 35076 100668
rect 35076 100612 35080 100668
rect 35016 100608 35080 100612
rect 35096 100668 35160 100672
rect 35096 100612 35100 100668
rect 35100 100612 35156 100668
rect 35156 100612 35160 100668
rect 35096 100608 35160 100612
rect 35176 100668 35240 100672
rect 35176 100612 35180 100668
rect 35180 100612 35236 100668
rect 35236 100612 35240 100668
rect 35176 100608 35240 100612
rect 65656 100668 65720 100672
rect 65656 100612 65660 100668
rect 65660 100612 65716 100668
rect 65716 100612 65720 100668
rect 65656 100608 65720 100612
rect 65736 100668 65800 100672
rect 65736 100612 65740 100668
rect 65740 100612 65796 100668
rect 65796 100612 65800 100668
rect 65736 100608 65800 100612
rect 65816 100668 65880 100672
rect 65816 100612 65820 100668
rect 65820 100612 65876 100668
rect 65876 100612 65880 100668
rect 65816 100608 65880 100612
rect 65896 100668 65960 100672
rect 65896 100612 65900 100668
rect 65900 100612 65956 100668
rect 65956 100612 65960 100668
rect 65896 100608 65960 100612
rect 19576 100124 19640 100128
rect 19576 100068 19580 100124
rect 19580 100068 19636 100124
rect 19636 100068 19640 100124
rect 19576 100064 19640 100068
rect 19656 100124 19720 100128
rect 19656 100068 19660 100124
rect 19660 100068 19716 100124
rect 19716 100068 19720 100124
rect 19656 100064 19720 100068
rect 19736 100124 19800 100128
rect 19736 100068 19740 100124
rect 19740 100068 19796 100124
rect 19796 100068 19800 100124
rect 19736 100064 19800 100068
rect 19816 100124 19880 100128
rect 19816 100068 19820 100124
rect 19820 100068 19876 100124
rect 19876 100068 19880 100124
rect 19816 100064 19880 100068
rect 50296 100124 50360 100128
rect 50296 100068 50300 100124
rect 50300 100068 50356 100124
rect 50356 100068 50360 100124
rect 50296 100064 50360 100068
rect 50376 100124 50440 100128
rect 50376 100068 50380 100124
rect 50380 100068 50436 100124
rect 50436 100068 50440 100124
rect 50376 100064 50440 100068
rect 50456 100124 50520 100128
rect 50456 100068 50460 100124
rect 50460 100068 50516 100124
rect 50516 100068 50520 100124
rect 50456 100064 50520 100068
rect 50536 100124 50600 100128
rect 50536 100068 50540 100124
rect 50540 100068 50596 100124
rect 50596 100068 50600 100124
rect 50536 100064 50600 100068
rect 4216 99580 4280 99584
rect 4216 99524 4220 99580
rect 4220 99524 4276 99580
rect 4276 99524 4280 99580
rect 4216 99520 4280 99524
rect 4296 99580 4360 99584
rect 4296 99524 4300 99580
rect 4300 99524 4356 99580
rect 4356 99524 4360 99580
rect 4296 99520 4360 99524
rect 4376 99580 4440 99584
rect 4376 99524 4380 99580
rect 4380 99524 4436 99580
rect 4436 99524 4440 99580
rect 4376 99520 4440 99524
rect 4456 99580 4520 99584
rect 4456 99524 4460 99580
rect 4460 99524 4516 99580
rect 4516 99524 4520 99580
rect 4456 99520 4520 99524
rect 34936 99580 35000 99584
rect 34936 99524 34940 99580
rect 34940 99524 34996 99580
rect 34996 99524 35000 99580
rect 34936 99520 35000 99524
rect 35016 99580 35080 99584
rect 35016 99524 35020 99580
rect 35020 99524 35076 99580
rect 35076 99524 35080 99580
rect 35016 99520 35080 99524
rect 35096 99580 35160 99584
rect 35096 99524 35100 99580
rect 35100 99524 35156 99580
rect 35156 99524 35160 99580
rect 35096 99520 35160 99524
rect 35176 99580 35240 99584
rect 35176 99524 35180 99580
rect 35180 99524 35236 99580
rect 35236 99524 35240 99580
rect 35176 99520 35240 99524
rect 65656 99580 65720 99584
rect 65656 99524 65660 99580
rect 65660 99524 65716 99580
rect 65716 99524 65720 99580
rect 65656 99520 65720 99524
rect 65736 99580 65800 99584
rect 65736 99524 65740 99580
rect 65740 99524 65796 99580
rect 65796 99524 65800 99580
rect 65736 99520 65800 99524
rect 65816 99580 65880 99584
rect 65816 99524 65820 99580
rect 65820 99524 65876 99580
rect 65876 99524 65880 99580
rect 65816 99520 65880 99524
rect 65896 99580 65960 99584
rect 65896 99524 65900 99580
rect 65900 99524 65956 99580
rect 65956 99524 65960 99580
rect 65896 99520 65960 99524
rect 19576 99036 19640 99040
rect 19576 98980 19580 99036
rect 19580 98980 19636 99036
rect 19636 98980 19640 99036
rect 19576 98976 19640 98980
rect 19656 99036 19720 99040
rect 19656 98980 19660 99036
rect 19660 98980 19716 99036
rect 19716 98980 19720 99036
rect 19656 98976 19720 98980
rect 19736 99036 19800 99040
rect 19736 98980 19740 99036
rect 19740 98980 19796 99036
rect 19796 98980 19800 99036
rect 19736 98976 19800 98980
rect 19816 99036 19880 99040
rect 19816 98980 19820 99036
rect 19820 98980 19876 99036
rect 19876 98980 19880 99036
rect 19816 98976 19880 98980
rect 50296 99036 50360 99040
rect 50296 98980 50300 99036
rect 50300 98980 50356 99036
rect 50356 98980 50360 99036
rect 50296 98976 50360 98980
rect 50376 99036 50440 99040
rect 50376 98980 50380 99036
rect 50380 98980 50436 99036
rect 50436 98980 50440 99036
rect 50376 98976 50440 98980
rect 50456 99036 50520 99040
rect 50456 98980 50460 99036
rect 50460 98980 50516 99036
rect 50516 98980 50520 99036
rect 50456 98976 50520 98980
rect 50536 99036 50600 99040
rect 50536 98980 50540 99036
rect 50540 98980 50596 99036
rect 50596 98980 50600 99036
rect 50536 98976 50600 98980
rect 4216 98492 4280 98496
rect 4216 98436 4220 98492
rect 4220 98436 4276 98492
rect 4276 98436 4280 98492
rect 4216 98432 4280 98436
rect 4296 98492 4360 98496
rect 4296 98436 4300 98492
rect 4300 98436 4356 98492
rect 4356 98436 4360 98492
rect 4296 98432 4360 98436
rect 4376 98492 4440 98496
rect 4376 98436 4380 98492
rect 4380 98436 4436 98492
rect 4436 98436 4440 98492
rect 4376 98432 4440 98436
rect 4456 98492 4520 98496
rect 4456 98436 4460 98492
rect 4460 98436 4516 98492
rect 4516 98436 4520 98492
rect 4456 98432 4520 98436
rect 34936 98492 35000 98496
rect 34936 98436 34940 98492
rect 34940 98436 34996 98492
rect 34996 98436 35000 98492
rect 34936 98432 35000 98436
rect 35016 98492 35080 98496
rect 35016 98436 35020 98492
rect 35020 98436 35076 98492
rect 35076 98436 35080 98492
rect 35016 98432 35080 98436
rect 35096 98492 35160 98496
rect 35096 98436 35100 98492
rect 35100 98436 35156 98492
rect 35156 98436 35160 98492
rect 35096 98432 35160 98436
rect 35176 98492 35240 98496
rect 35176 98436 35180 98492
rect 35180 98436 35236 98492
rect 35236 98436 35240 98492
rect 35176 98432 35240 98436
rect 65656 98492 65720 98496
rect 65656 98436 65660 98492
rect 65660 98436 65716 98492
rect 65716 98436 65720 98492
rect 65656 98432 65720 98436
rect 65736 98492 65800 98496
rect 65736 98436 65740 98492
rect 65740 98436 65796 98492
rect 65796 98436 65800 98492
rect 65736 98432 65800 98436
rect 65816 98492 65880 98496
rect 65816 98436 65820 98492
rect 65820 98436 65876 98492
rect 65876 98436 65880 98492
rect 65816 98432 65880 98436
rect 65896 98492 65960 98496
rect 65896 98436 65900 98492
rect 65900 98436 65956 98492
rect 65956 98436 65960 98492
rect 65896 98432 65960 98436
rect 19576 97948 19640 97952
rect 19576 97892 19580 97948
rect 19580 97892 19636 97948
rect 19636 97892 19640 97948
rect 19576 97888 19640 97892
rect 19656 97948 19720 97952
rect 19656 97892 19660 97948
rect 19660 97892 19716 97948
rect 19716 97892 19720 97948
rect 19656 97888 19720 97892
rect 19736 97948 19800 97952
rect 19736 97892 19740 97948
rect 19740 97892 19796 97948
rect 19796 97892 19800 97948
rect 19736 97888 19800 97892
rect 19816 97948 19880 97952
rect 19816 97892 19820 97948
rect 19820 97892 19876 97948
rect 19876 97892 19880 97948
rect 19816 97888 19880 97892
rect 50296 97948 50360 97952
rect 50296 97892 50300 97948
rect 50300 97892 50356 97948
rect 50356 97892 50360 97948
rect 50296 97888 50360 97892
rect 50376 97948 50440 97952
rect 50376 97892 50380 97948
rect 50380 97892 50436 97948
rect 50436 97892 50440 97948
rect 50376 97888 50440 97892
rect 50456 97948 50520 97952
rect 50456 97892 50460 97948
rect 50460 97892 50516 97948
rect 50516 97892 50520 97948
rect 50456 97888 50520 97892
rect 50536 97948 50600 97952
rect 50536 97892 50540 97948
rect 50540 97892 50596 97948
rect 50596 97892 50600 97948
rect 50536 97888 50600 97892
rect 4216 97404 4280 97408
rect 4216 97348 4220 97404
rect 4220 97348 4276 97404
rect 4276 97348 4280 97404
rect 4216 97344 4280 97348
rect 4296 97404 4360 97408
rect 4296 97348 4300 97404
rect 4300 97348 4356 97404
rect 4356 97348 4360 97404
rect 4296 97344 4360 97348
rect 4376 97404 4440 97408
rect 4376 97348 4380 97404
rect 4380 97348 4436 97404
rect 4436 97348 4440 97404
rect 4376 97344 4440 97348
rect 4456 97404 4520 97408
rect 4456 97348 4460 97404
rect 4460 97348 4516 97404
rect 4516 97348 4520 97404
rect 4456 97344 4520 97348
rect 34936 97404 35000 97408
rect 34936 97348 34940 97404
rect 34940 97348 34996 97404
rect 34996 97348 35000 97404
rect 34936 97344 35000 97348
rect 35016 97404 35080 97408
rect 35016 97348 35020 97404
rect 35020 97348 35076 97404
rect 35076 97348 35080 97404
rect 35016 97344 35080 97348
rect 35096 97404 35160 97408
rect 35096 97348 35100 97404
rect 35100 97348 35156 97404
rect 35156 97348 35160 97404
rect 35096 97344 35160 97348
rect 35176 97404 35240 97408
rect 35176 97348 35180 97404
rect 35180 97348 35236 97404
rect 35236 97348 35240 97404
rect 35176 97344 35240 97348
rect 65656 97404 65720 97408
rect 65656 97348 65660 97404
rect 65660 97348 65716 97404
rect 65716 97348 65720 97404
rect 65656 97344 65720 97348
rect 65736 97404 65800 97408
rect 65736 97348 65740 97404
rect 65740 97348 65796 97404
rect 65796 97348 65800 97404
rect 65736 97344 65800 97348
rect 65816 97404 65880 97408
rect 65816 97348 65820 97404
rect 65820 97348 65876 97404
rect 65876 97348 65880 97404
rect 65816 97344 65880 97348
rect 65896 97404 65960 97408
rect 65896 97348 65900 97404
rect 65900 97348 65956 97404
rect 65956 97348 65960 97404
rect 65896 97344 65960 97348
rect 19576 96860 19640 96864
rect 19576 96804 19580 96860
rect 19580 96804 19636 96860
rect 19636 96804 19640 96860
rect 19576 96800 19640 96804
rect 19656 96860 19720 96864
rect 19656 96804 19660 96860
rect 19660 96804 19716 96860
rect 19716 96804 19720 96860
rect 19656 96800 19720 96804
rect 19736 96860 19800 96864
rect 19736 96804 19740 96860
rect 19740 96804 19796 96860
rect 19796 96804 19800 96860
rect 19736 96800 19800 96804
rect 19816 96860 19880 96864
rect 19816 96804 19820 96860
rect 19820 96804 19876 96860
rect 19876 96804 19880 96860
rect 19816 96800 19880 96804
rect 50296 96860 50360 96864
rect 50296 96804 50300 96860
rect 50300 96804 50356 96860
rect 50356 96804 50360 96860
rect 50296 96800 50360 96804
rect 50376 96860 50440 96864
rect 50376 96804 50380 96860
rect 50380 96804 50436 96860
rect 50436 96804 50440 96860
rect 50376 96800 50440 96804
rect 50456 96860 50520 96864
rect 50456 96804 50460 96860
rect 50460 96804 50516 96860
rect 50516 96804 50520 96860
rect 50456 96800 50520 96804
rect 50536 96860 50600 96864
rect 50536 96804 50540 96860
rect 50540 96804 50596 96860
rect 50596 96804 50600 96860
rect 50536 96800 50600 96804
rect 4216 96316 4280 96320
rect 4216 96260 4220 96316
rect 4220 96260 4276 96316
rect 4276 96260 4280 96316
rect 4216 96256 4280 96260
rect 4296 96316 4360 96320
rect 4296 96260 4300 96316
rect 4300 96260 4356 96316
rect 4356 96260 4360 96316
rect 4296 96256 4360 96260
rect 4376 96316 4440 96320
rect 4376 96260 4380 96316
rect 4380 96260 4436 96316
rect 4436 96260 4440 96316
rect 4376 96256 4440 96260
rect 4456 96316 4520 96320
rect 4456 96260 4460 96316
rect 4460 96260 4516 96316
rect 4516 96260 4520 96316
rect 4456 96256 4520 96260
rect 34936 96316 35000 96320
rect 34936 96260 34940 96316
rect 34940 96260 34996 96316
rect 34996 96260 35000 96316
rect 34936 96256 35000 96260
rect 35016 96316 35080 96320
rect 35016 96260 35020 96316
rect 35020 96260 35076 96316
rect 35076 96260 35080 96316
rect 35016 96256 35080 96260
rect 35096 96316 35160 96320
rect 35096 96260 35100 96316
rect 35100 96260 35156 96316
rect 35156 96260 35160 96316
rect 35096 96256 35160 96260
rect 35176 96316 35240 96320
rect 35176 96260 35180 96316
rect 35180 96260 35236 96316
rect 35236 96260 35240 96316
rect 35176 96256 35240 96260
rect 65656 96316 65720 96320
rect 65656 96260 65660 96316
rect 65660 96260 65716 96316
rect 65716 96260 65720 96316
rect 65656 96256 65720 96260
rect 65736 96316 65800 96320
rect 65736 96260 65740 96316
rect 65740 96260 65796 96316
rect 65796 96260 65800 96316
rect 65736 96256 65800 96260
rect 65816 96316 65880 96320
rect 65816 96260 65820 96316
rect 65820 96260 65876 96316
rect 65876 96260 65880 96316
rect 65816 96256 65880 96260
rect 65896 96316 65960 96320
rect 65896 96260 65900 96316
rect 65900 96260 65956 96316
rect 65956 96260 65960 96316
rect 65896 96256 65960 96260
rect 19576 95772 19640 95776
rect 19576 95716 19580 95772
rect 19580 95716 19636 95772
rect 19636 95716 19640 95772
rect 19576 95712 19640 95716
rect 19656 95772 19720 95776
rect 19656 95716 19660 95772
rect 19660 95716 19716 95772
rect 19716 95716 19720 95772
rect 19656 95712 19720 95716
rect 19736 95772 19800 95776
rect 19736 95716 19740 95772
rect 19740 95716 19796 95772
rect 19796 95716 19800 95772
rect 19736 95712 19800 95716
rect 19816 95772 19880 95776
rect 19816 95716 19820 95772
rect 19820 95716 19876 95772
rect 19876 95716 19880 95772
rect 19816 95712 19880 95716
rect 50296 95772 50360 95776
rect 50296 95716 50300 95772
rect 50300 95716 50356 95772
rect 50356 95716 50360 95772
rect 50296 95712 50360 95716
rect 50376 95772 50440 95776
rect 50376 95716 50380 95772
rect 50380 95716 50436 95772
rect 50436 95716 50440 95772
rect 50376 95712 50440 95716
rect 50456 95772 50520 95776
rect 50456 95716 50460 95772
rect 50460 95716 50516 95772
rect 50516 95716 50520 95772
rect 50456 95712 50520 95716
rect 50536 95772 50600 95776
rect 50536 95716 50540 95772
rect 50540 95716 50596 95772
rect 50596 95716 50600 95772
rect 50536 95712 50600 95716
rect 4216 95228 4280 95232
rect 4216 95172 4220 95228
rect 4220 95172 4276 95228
rect 4276 95172 4280 95228
rect 4216 95168 4280 95172
rect 4296 95228 4360 95232
rect 4296 95172 4300 95228
rect 4300 95172 4356 95228
rect 4356 95172 4360 95228
rect 4296 95168 4360 95172
rect 4376 95228 4440 95232
rect 4376 95172 4380 95228
rect 4380 95172 4436 95228
rect 4436 95172 4440 95228
rect 4376 95168 4440 95172
rect 4456 95228 4520 95232
rect 4456 95172 4460 95228
rect 4460 95172 4516 95228
rect 4516 95172 4520 95228
rect 4456 95168 4520 95172
rect 34936 95228 35000 95232
rect 34936 95172 34940 95228
rect 34940 95172 34996 95228
rect 34996 95172 35000 95228
rect 34936 95168 35000 95172
rect 35016 95228 35080 95232
rect 35016 95172 35020 95228
rect 35020 95172 35076 95228
rect 35076 95172 35080 95228
rect 35016 95168 35080 95172
rect 35096 95228 35160 95232
rect 35096 95172 35100 95228
rect 35100 95172 35156 95228
rect 35156 95172 35160 95228
rect 35096 95168 35160 95172
rect 35176 95228 35240 95232
rect 35176 95172 35180 95228
rect 35180 95172 35236 95228
rect 35236 95172 35240 95228
rect 35176 95168 35240 95172
rect 65656 95228 65720 95232
rect 65656 95172 65660 95228
rect 65660 95172 65716 95228
rect 65716 95172 65720 95228
rect 65656 95168 65720 95172
rect 65736 95228 65800 95232
rect 65736 95172 65740 95228
rect 65740 95172 65796 95228
rect 65796 95172 65800 95228
rect 65736 95168 65800 95172
rect 65816 95228 65880 95232
rect 65816 95172 65820 95228
rect 65820 95172 65876 95228
rect 65876 95172 65880 95228
rect 65816 95168 65880 95172
rect 65896 95228 65960 95232
rect 65896 95172 65900 95228
rect 65900 95172 65956 95228
rect 65956 95172 65960 95228
rect 65896 95168 65960 95172
rect 19576 94684 19640 94688
rect 19576 94628 19580 94684
rect 19580 94628 19636 94684
rect 19636 94628 19640 94684
rect 19576 94624 19640 94628
rect 19656 94684 19720 94688
rect 19656 94628 19660 94684
rect 19660 94628 19716 94684
rect 19716 94628 19720 94684
rect 19656 94624 19720 94628
rect 19736 94684 19800 94688
rect 19736 94628 19740 94684
rect 19740 94628 19796 94684
rect 19796 94628 19800 94684
rect 19736 94624 19800 94628
rect 19816 94684 19880 94688
rect 19816 94628 19820 94684
rect 19820 94628 19876 94684
rect 19876 94628 19880 94684
rect 19816 94624 19880 94628
rect 50296 94684 50360 94688
rect 50296 94628 50300 94684
rect 50300 94628 50356 94684
rect 50356 94628 50360 94684
rect 50296 94624 50360 94628
rect 50376 94684 50440 94688
rect 50376 94628 50380 94684
rect 50380 94628 50436 94684
rect 50436 94628 50440 94684
rect 50376 94624 50440 94628
rect 50456 94684 50520 94688
rect 50456 94628 50460 94684
rect 50460 94628 50516 94684
rect 50516 94628 50520 94684
rect 50456 94624 50520 94628
rect 50536 94684 50600 94688
rect 50536 94628 50540 94684
rect 50540 94628 50596 94684
rect 50596 94628 50600 94684
rect 50536 94624 50600 94628
rect 4216 94140 4280 94144
rect 4216 94084 4220 94140
rect 4220 94084 4276 94140
rect 4276 94084 4280 94140
rect 4216 94080 4280 94084
rect 4296 94140 4360 94144
rect 4296 94084 4300 94140
rect 4300 94084 4356 94140
rect 4356 94084 4360 94140
rect 4296 94080 4360 94084
rect 4376 94140 4440 94144
rect 4376 94084 4380 94140
rect 4380 94084 4436 94140
rect 4436 94084 4440 94140
rect 4376 94080 4440 94084
rect 4456 94140 4520 94144
rect 4456 94084 4460 94140
rect 4460 94084 4516 94140
rect 4516 94084 4520 94140
rect 4456 94080 4520 94084
rect 34936 94140 35000 94144
rect 34936 94084 34940 94140
rect 34940 94084 34996 94140
rect 34996 94084 35000 94140
rect 34936 94080 35000 94084
rect 35016 94140 35080 94144
rect 35016 94084 35020 94140
rect 35020 94084 35076 94140
rect 35076 94084 35080 94140
rect 35016 94080 35080 94084
rect 35096 94140 35160 94144
rect 35096 94084 35100 94140
rect 35100 94084 35156 94140
rect 35156 94084 35160 94140
rect 35096 94080 35160 94084
rect 35176 94140 35240 94144
rect 35176 94084 35180 94140
rect 35180 94084 35236 94140
rect 35236 94084 35240 94140
rect 35176 94080 35240 94084
rect 65656 94140 65720 94144
rect 65656 94084 65660 94140
rect 65660 94084 65716 94140
rect 65716 94084 65720 94140
rect 65656 94080 65720 94084
rect 65736 94140 65800 94144
rect 65736 94084 65740 94140
rect 65740 94084 65796 94140
rect 65796 94084 65800 94140
rect 65736 94080 65800 94084
rect 65816 94140 65880 94144
rect 65816 94084 65820 94140
rect 65820 94084 65876 94140
rect 65876 94084 65880 94140
rect 65816 94080 65880 94084
rect 65896 94140 65960 94144
rect 65896 94084 65900 94140
rect 65900 94084 65956 94140
rect 65956 94084 65960 94140
rect 65896 94080 65960 94084
rect 19576 93596 19640 93600
rect 19576 93540 19580 93596
rect 19580 93540 19636 93596
rect 19636 93540 19640 93596
rect 19576 93536 19640 93540
rect 19656 93596 19720 93600
rect 19656 93540 19660 93596
rect 19660 93540 19716 93596
rect 19716 93540 19720 93596
rect 19656 93536 19720 93540
rect 19736 93596 19800 93600
rect 19736 93540 19740 93596
rect 19740 93540 19796 93596
rect 19796 93540 19800 93596
rect 19736 93536 19800 93540
rect 19816 93596 19880 93600
rect 19816 93540 19820 93596
rect 19820 93540 19876 93596
rect 19876 93540 19880 93596
rect 19816 93536 19880 93540
rect 50296 93596 50360 93600
rect 50296 93540 50300 93596
rect 50300 93540 50356 93596
rect 50356 93540 50360 93596
rect 50296 93536 50360 93540
rect 50376 93596 50440 93600
rect 50376 93540 50380 93596
rect 50380 93540 50436 93596
rect 50436 93540 50440 93596
rect 50376 93536 50440 93540
rect 50456 93596 50520 93600
rect 50456 93540 50460 93596
rect 50460 93540 50516 93596
rect 50516 93540 50520 93596
rect 50456 93536 50520 93540
rect 50536 93596 50600 93600
rect 50536 93540 50540 93596
rect 50540 93540 50596 93596
rect 50596 93540 50600 93596
rect 50536 93536 50600 93540
rect 4216 93052 4280 93056
rect 4216 92996 4220 93052
rect 4220 92996 4276 93052
rect 4276 92996 4280 93052
rect 4216 92992 4280 92996
rect 4296 93052 4360 93056
rect 4296 92996 4300 93052
rect 4300 92996 4356 93052
rect 4356 92996 4360 93052
rect 4296 92992 4360 92996
rect 4376 93052 4440 93056
rect 4376 92996 4380 93052
rect 4380 92996 4436 93052
rect 4436 92996 4440 93052
rect 4376 92992 4440 92996
rect 4456 93052 4520 93056
rect 4456 92996 4460 93052
rect 4460 92996 4516 93052
rect 4516 92996 4520 93052
rect 4456 92992 4520 92996
rect 34936 93052 35000 93056
rect 34936 92996 34940 93052
rect 34940 92996 34996 93052
rect 34996 92996 35000 93052
rect 34936 92992 35000 92996
rect 35016 93052 35080 93056
rect 35016 92996 35020 93052
rect 35020 92996 35076 93052
rect 35076 92996 35080 93052
rect 35016 92992 35080 92996
rect 35096 93052 35160 93056
rect 35096 92996 35100 93052
rect 35100 92996 35156 93052
rect 35156 92996 35160 93052
rect 35096 92992 35160 92996
rect 35176 93052 35240 93056
rect 35176 92996 35180 93052
rect 35180 92996 35236 93052
rect 35236 92996 35240 93052
rect 35176 92992 35240 92996
rect 65656 93052 65720 93056
rect 65656 92996 65660 93052
rect 65660 92996 65716 93052
rect 65716 92996 65720 93052
rect 65656 92992 65720 92996
rect 65736 93052 65800 93056
rect 65736 92996 65740 93052
rect 65740 92996 65796 93052
rect 65796 92996 65800 93052
rect 65736 92992 65800 92996
rect 65816 93052 65880 93056
rect 65816 92996 65820 93052
rect 65820 92996 65876 93052
rect 65876 92996 65880 93052
rect 65816 92992 65880 92996
rect 65896 93052 65960 93056
rect 65896 92996 65900 93052
rect 65900 92996 65956 93052
rect 65956 92996 65960 93052
rect 65896 92992 65960 92996
rect 19576 92508 19640 92512
rect 19576 92452 19580 92508
rect 19580 92452 19636 92508
rect 19636 92452 19640 92508
rect 19576 92448 19640 92452
rect 19656 92508 19720 92512
rect 19656 92452 19660 92508
rect 19660 92452 19716 92508
rect 19716 92452 19720 92508
rect 19656 92448 19720 92452
rect 19736 92508 19800 92512
rect 19736 92452 19740 92508
rect 19740 92452 19796 92508
rect 19796 92452 19800 92508
rect 19736 92448 19800 92452
rect 19816 92508 19880 92512
rect 19816 92452 19820 92508
rect 19820 92452 19876 92508
rect 19876 92452 19880 92508
rect 19816 92448 19880 92452
rect 50296 92508 50360 92512
rect 50296 92452 50300 92508
rect 50300 92452 50356 92508
rect 50356 92452 50360 92508
rect 50296 92448 50360 92452
rect 50376 92508 50440 92512
rect 50376 92452 50380 92508
rect 50380 92452 50436 92508
rect 50436 92452 50440 92508
rect 50376 92448 50440 92452
rect 50456 92508 50520 92512
rect 50456 92452 50460 92508
rect 50460 92452 50516 92508
rect 50516 92452 50520 92508
rect 50456 92448 50520 92452
rect 50536 92508 50600 92512
rect 50536 92452 50540 92508
rect 50540 92452 50596 92508
rect 50596 92452 50600 92508
rect 50536 92448 50600 92452
rect 4216 91964 4280 91968
rect 4216 91908 4220 91964
rect 4220 91908 4276 91964
rect 4276 91908 4280 91964
rect 4216 91904 4280 91908
rect 4296 91964 4360 91968
rect 4296 91908 4300 91964
rect 4300 91908 4356 91964
rect 4356 91908 4360 91964
rect 4296 91904 4360 91908
rect 4376 91964 4440 91968
rect 4376 91908 4380 91964
rect 4380 91908 4436 91964
rect 4436 91908 4440 91964
rect 4376 91904 4440 91908
rect 4456 91964 4520 91968
rect 4456 91908 4460 91964
rect 4460 91908 4516 91964
rect 4516 91908 4520 91964
rect 4456 91904 4520 91908
rect 34936 91964 35000 91968
rect 34936 91908 34940 91964
rect 34940 91908 34996 91964
rect 34996 91908 35000 91964
rect 34936 91904 35000 91908
rect 35016 91964 35080 91968
rect 35016 91908 35020 91964
rect 35020 91908 35076 91964
rect 35076 91908 35080 91964
rect 35016 91904 35080 91908
rect 35096 91964 35160 91968
rect 35096 91908 35100 91964
rect 35100 91908 35156 91964
rect 35156 91908 35160 91964
rect 35096 91904 35160 91908
rect 35176 91964 35240 91968
rect 35176 91908 35180 91964
rect 35180 91908 35236 91964
rect 35236 91908 35240 91964
rect 35176 91904 35240 91908
rect 65656 91964 65720 91968
rect 65656 91908 65660 91964
rect 65660 91908 65716 91964
rect 65716 91908 65720 91964
rect 65656 91904 65720 91908
rect 65736 91964 65800 91968
rect 65736 91908 65740 91964
rect 65740 91908 65796 91964
rect 65796 91908 65800 91964
rect 65736 91904 65800 91908
rect 65816 91964 65880 91968
rect 65816 91908 65820 91964
rect 65820 91908 65876 91964
rect 65876 91908 65880 91964
rect 65816 91904 65880 91908
rect 65896 91964 65960 91968
rect 65896 91908 65900 91964
rect 65900 91908 65956 91964
rect 65956 91908 65960 91964
rect 65896 91904 65960 91908
rect 19576 91420 19640 91424
rect 19576 91364 19580 91420
rect 19580 91364 19636 91420
rect 19636 91364 19640 91420
rect 19576 91360 19640 91364
rect 19656 91420 19720 91424
rect 19656 91364 19660 91420
rect 19660 91364 19716 91420
rect 19716 91364 19720 91420
rect 19656 91360 19720 91364
rect 19736 91420 19800 91424
rect 19736 91364 19740 91420
rect 19740 91364 19796 91420
rect 19796 91364 19800 91420
rect 19736 91360 19800 91364
rect 19816 91420 19880 91424
rect 19816 91364 19820 91420
rect 19820 91364 19876 91420
rect 19876 91364 19880 91420
rect 19816 91360 19880 91364
rect 50296 91420 50360 91424
rect 50296 91364 50300 91420
rect 50300 91364 50356 91420
rect 50356 91364 50360 91420
rect 50296 91360 50360 91364
rect 50376 91420 50440 91424
rect 50376 91364 50380 91420
rect 50380 91364 50436 91420
rect 50436 91364 50440 91420
rect 50376 91360 50440 91364
rect 50456 91420 50520 91424
rect 50456 91364 50460 91420
rect 50460 91364 50516 91420
rect 50516 91364 50520 91420
rect 50456 91360 50520 91364
rect 50536 91420 50600 91424
rect 50536 91364 50540 91420
rect 50540 91364 50596 91420
rect 50596 91364 50600 91420
rect 50536 91360 50600 91364
rect 4216 90876 4280 90880
rect 4216 90820 4220 90876
rect 4220 90820 4276 90876
rect 4276 90820 4280 90876
rect 4216 90816 4280 90820
rect 4296 90876 4360 90880
rect 4296 90820 4300 90876
rect 4300 90820 4356 90876
rect 4356 90820 4360 90876
rect 4296 90816 4360 90820
rect 4376 90876 4440 90880
rect 4376 90820 4380 90876
rect 4380 90820 4436 90876
rect 4436 90820 4440 90876
rect 4376 90816 4440 90820
rect 4456 90876 4520 90880
rect 4456 90820 4460 90876
rect 4460 90820 4516 90876
rect 4516 90820 4520 90876
rect 4456 90816 4520 90820
rect 34936 90876 35000 90880
rect 34936 90820 34940 90876
rect 34940 90820 34996 90876
rect 34996 90820 35000 90876
rect 34936 90816 35000 90820
rect 35016 90876 35080 90880
rect 35016 90820 35020 90876
rect 35020 90820 35076 90876
rect 35076 90820 35080 90876
rect 35016 90816 35080 90820
rect 35096 90876 35160 90880
rect 35096 90820 35100 90876
rect 35100 90820 35156 90876
rect 35156 90820 35160 90876
rect 35096 90816 35160 90820
rect 35176 90876 35240 90880
rect 35176 90820 35180 90876
rect 35180 90820 35236 90876
rect 35236 90820 35240 90876
rect 35176 90816 35240 90820
rect 65656 90876 65720 90880
rect 65656 90820 65660 90876
rect 65660 90820 65716 90876
rect 65716 90820 65720 90876
rect 65656 90816 65720 90820
rect 65736 90876 65800 90880
rect 65736 90820 65740 90876
rect 65740 90820 65796 90876
rect 65796 90820 65800 90876
rect 65736 90816 65800 90820
rect 65816 90876 65880 90880
rect 65816 90820 65820 90876
rect 65820 90820 65876 90876
rect 65876 90820 65880 90876
rect 65816 90816 65880 90820
rect 65896 90876 65960 90880
rect 65896 90820 65900 90876
rect 65900 90820 65956 90876
rect 65956 90820 65960 90876
rect 65896 90816 65960 90820
rect 19576 90332 19640 90336
rect 19576 90276 19580 90332
rect 19580 90276 19636 90332
rect 19636 90276 19640 90332
rect 19576 90272 19640 90276
rect 19656 90332 19720 90336
rect 19656 90276 19660 90332
rect 19660 90276 19716 90332
rect 19716 90276 19720 90332
rect 19656 90272 19720 90276
rect 19736 90332 19800 90336
rect 19736 90276 19740 90332
rect 19740 90276 19796 90332
rect 19796 90276 19800 90332
rect 19736 90272 19800 90276
rect 19816 90332 19880 90336
rect 19816 90276 19820 90332
rect 19820 90276 19876 90332
rect 19876 90276 19880 90332
rect 19816 90272 19880 90276
rect 50296 90332 50360 90336
rect 50296 90276 50300 90332
rect 50300 90276 50356 90332
rect 50356 90276 50360 90332
rect 50296 90272 50360 90276
rect 50376 90332 50440 90336
rect 50376 90276 50380 90332
rect 50380 90276 50436 90332
rect 50436 90276 50440 90332
rect 50376 90272 50440 90276
rect 50456 90332 50520 90336
rect 50456 90276 50460 90332
rect 50460 90276 50516 90332
rect 50516 90276 50520 90332
rect 50456 90272 50520 90276
rect 50536 90332 50600 90336
rect 50536 90276 50540 90332
rect 50540 90276 50596 90332
rect 50596 90276 50600 90332
rect 50536 90272 50600 90276
rect 4216 89788 4280 89792
rect 4216 89732 4220 89788
rect 4220 89732 4276 89788
rect 4276 89732 4280 89788
rect 4216 89728 4280 89732
rect 4296 89788 4360 89792
rect 4296 89732 4300 89788
rect 4300 89732 4356 89788
rect 4356 89732 4360 89788
rect 4296 89728 4360 89732
rect 4376 89788 4440 89792
rect 4376 89732 4380 89788
rect 4380 89732 4436 89788
rect 4436 89732 4440 89788
rect 4376 89728 4440 89732
rect 4456 89788 4520 89792
rect 4456 89732 4460 89788
rect 4460 89732 4516 89788
rect 4516 89732 4520 89788
rect 4456 89728 4520 89732
rect 34936 89788 35000 89792
rect 34936 89732 34940 89788
rect 34940 89732 34996 89788
rect 34996 89732 35000 89788
rect 34936 89728 35000 89732
rect 35016 89788 35080 89792
rect 35016 89732 35020 89788
rect 35020 89732 35076 89788
rect 35076 89732 35080 89788
rect 35016 89728 35080 89732
rect 35096 89788 35160 89792
rect 35096 89732 35100 89788
rect 35100 89732 35156 89788
rect 35156 89732 35160 89788
rect 35096 89728 35160 89732
rect 35176 89788 35240 89792
rect 35176 89732 35180 89788
rect 35180 89732 35236 89788
rect 35236 89732 35240 89788
rect 35176 89728 35240 89732
rect 65656 89788 65720 89792
rect 65656 89732 65660 89788
rect 65660 89732 65716 89788
rect 65716 89732 65720 89788
rect 65656 89728 65720 89732
rect 65736 89788 65800 89792
rect 65736 89732 65740 89788
rect 65740 89732 65796 89788
rect 65796 89732 65800 89788
rect 65736 89728 65800 89732
rect 65816 89788 65880 89792
rect 65816 89732 65820 89788
rect 65820 89732 65876 89788
rect 65876 89732 65880 89788
rect 65816 89728 65880 89732
rect 65896 89788 65960 89792
rect 65896 89732 65900 89788
rect 65900 89732 65956 89788
rect 65956 89732 65960 89788
rect 65896 89728 65960 89732
rect 19576 89244 19640 89248
rect 19576 89188 19580 89244
rect 19580 89188 19636 89244
rect 19636 89188 19640 89244
rect 19576 89184 19640 89188
rect 19656 89244 19720 89248
rect 19656 89188 19660 89244
rect 19660 89188 19716 89244
rect 19716 89188 19720 89244
rect 19656 89184 19720 89188
rect 19736 89244 19800 89248
rect 19736 89188 19740 89244
rect 19740 89188 19796 89244
rect 19796 89188 19800 89244
rect 19736 89184 19800 89188
rect 19816 89244 19880 89248
rect 19816 89188 19820 89244
rect 19820 89188 19876 89244
rect 19876 89188 19880 89244
rect 19816 89184 19880 89188
rect 50296 89244 50360 89248
rect 50296 89188 50300 89244
rect 50300 89188 50356 89244
rect 50356 89188 50360 89244
rect 50296 89184 50360 89188
rect 50376 89244 50440 89248
rect 50376 89188 50380 89244
rect 50380 89188 50436 89244
rect 50436 89188 50440 89244
rect 50376 89184 50440 89188
rect 50456 89244 50520 89248
rect 50456 89188 50460 89244
rect 50460 89188 50516 89244
rect 50516 89188 50520 89244
rect 50456 89184 50520 89188
rect 50536 89244 50600 89248
rect 50536 89188 50540 89244
rect 50540 89188 50596 89244
rect 50596 89188 50600 89244
rect 50536 89184 50600 89188
rect 4216 88700 4280 88704
rect 4216 88644 4220 88700
rect 4220 88644 4276 88700
rect 4276 88644 4280 88700
rect 4216 88640 4280 88644
rect 4296 88700 4360 88704
rect 4296 88644 4300 88700
rect 4300 88644 4356 88700
rect 4356 88644 4360 88700
rect 4296 88640 4360 88644
rect 4376 88700 4440 88704
rect 4376 88644 4380 88700
rect 4380 88644 4436 88700
rect 4436 88644 4440 88700
rect 4376 88640 4440 88644
rect 4456 88700 4520 88704
rect 4456 88644 4460 88700
rect 4460 88644 4516 88700
rect 4516 88644 4520 88700
rect 4456 88640 4520 88644
rect 34936 88700 35000 88704
rect 34936 88644 34940 88700
rect 34940 88644 34996 88700
rect 34996 88644 35000 88700
rect 34936 88640 35000 88644
rect 35016 88700 35080 88704
rect 35016 88644 35020 88700
rect 35020 88644 35076 88700
rect 35076 88644 35080 88700
rect 35016 88640 35080 88644
rect 35096 88700 35160 88704
rect 35096 88644 35100 88700
rect 35100 88644 35156 88700
rect 35156 88644 35160 88700
rect 35096 88640 35160 88644
rect 35176 88700 35240 88704
rect 35176 88644 35180 88700
rect 35180 88644 35236 88700
rect 35236 88644 35240 88700
rect 35176 88640 35240 88644
rect 65656 88700 65720 88704
rect 65656 88644 65660 88700
rect 65660 88644 65716 88700
rect 65716 88644 65720 88700
rect 65656 88640 65720 88644
rect 65736 88700 65800 88704
rect 65736 88644 65740 88700
rect 65740 88644 65796 88700
rect 65796 88644 65800 88700
rect 65736 88640 65800 88644
rect 65816 88700 65880 88704
rect 65816 88644 65820 88700
rect 65820 88644 65876 88700
rect 65876 88644 65880 88700
rect 65816 88640 65880 88644
rect 65896 88700 65960 88704
rect 65896 88644 65900 88700
rect 65900 88644 65956 88700
rect 65956 88644 65960 88700
rect 65896 88640 65960 88644
rect 19576 88156 19640 88160
rect 19576 88100 19580 88156
rect 19580 88100 19636 88156
rect 19636 88100 19640 88156
rect 19576 88096 19640 88100
rect 19656 88156 19720 88160
rect 19656 88100 19660 88156
rect 19660 88100 19716 88156
rect 19716 88100 19720 88156
rect 19656 88096 19720 88100
rect 19736 88156 19800 88160
rect 19736 88100 19740 88156
rect 19740 88100 19796 88156
rect 19796 88100 19800 88156
rect 19736 88096 19800 88100
rect 19816 88156 19880 88160
rect 19816 88100 19820 88156
rect 19820 88100 19876 88156
rect 19876 88100 19880 88156
rect 19816 88096 19880 88100
rect 50296 88156 50360 88160
rect 50296 88100 50300 88156
rect 50300 88100 50356 88156
rect 50356 88100 50360 88156
rect 50296 88096 50360 88100
rect 50376 88156 50440 88160
rect 50376 88100 50380 88156
rect 50380 88100 50436 88156
rect 50436 88100 50440 88156
rect 50376 88096 50440 88100
rect 50456 88156 50520 88160
rect 50456 88100 50460 88156
rect 50460 88100 50516 88156
rect 50516 88100 50520 88156
rect 50456 88096 50520 88100
rect 50536 88156 50600 88160
rect 50536 88100 50540 88156
rect 50540 88100 50596 88156
rect 50596 88100 50600 88156
rect 50536 88096 50600 88100
rect 4216 87612 4280 87616
rect 4216 87556 4220 87612
rect 4220 87556 4276 87612
rect 4276 87556 4280 87612
rect 4216 87552 4280 87556
rect 4296 87612 4360 87616
rect 4296 87556 4300 87612
rect 4300 87556 4356 87612
rect 4356 87556 4360 87612
rect 4296 87552 4360 87556
rect 4376 87612 4440 87616
rect 4376 87556 4380 87612
rect 4380 87556 4436 87612
rect 4436 87556 4440 87612
rect 4376 87552 4440 87556
rect 4456 87612 4520 87616
rect 4456 87556 4460 87612
rect 4460 87556 4516 87612
rect 4516 87556 4520 87612
rect 4456 87552 4520 87556
rect 34936 87612 35000 87616
rect 34936 87556 34940 87612
rect 34940 87556 34996 87612
rect 34996 87556 35000 87612
rect 34936 87552 35000 87556
rect 35016 87612 35080 87616
rect 35016 87556 35020 87612
rect 35020 87556 35076 87612
rect 35076 87556 35080 87612
rect 35016 87552 35080 87556
rect 35096 87612 35160 87616
rect 35096 87556 35100 87612
rect 35100 87556 35156 87612
rect 35156 87556 35160 87612
rect 35096 87552 35160 87556
rect 35176 87612 35240 87616
rect 35176 87556 35180 87612
rect 35180 87556 35236 87612
rect 35236 87556 35240 87612
rect 35176 87552 35240 87556
rect 65656 87612 65720 87616
rect 65656 87556 65660 87612
rect 65660 87556 65716 87612
rect 65716 87556 65720 87612
rect 65656 87552 65720 87556
rect 65736 87612 65800 87616
rect 65736 87556 65740 87612
rect 65740 87556 65796 87612
rect 65796 87556 65800 87612
rect 65736 87552 65800 87556
rect 65816 87612 65880 87616
rect 65816 87556 65820 87612
rect 65820 87556 65876 87612
rect 65876 87556 65880 87612
rect 65816 87552 65880 87556
rect 65896 87612 65960 87616
rect 65896 87556 65900 87612
rect 65900 87556 65956 87612
rect 65956 87556 65960 87612
rect 65896 87552 65960 87556
rect 19576 87068 19640 87072
rect 19576 87012 19580 87068
rect 19580 87012 19636 87068
rect 19636 87012 19640 87068
rect 19576 87008 19640 87012
rect 19656 87068 19720 87072
rect 19656 87012 19660 87068
rect 19660 87012 19716 87068
rect 19716 87012 19720 87068
rect 19656 87008 19720 87012
rect 19736 87068 19800 87072
rect 19736 87012 19740 87068
rect 19740 87012 19796 87068
rect 19796 87012 19800 87068
rect 19736 87008 19800 87012
rect 19816 87068 19880 87072
rect 19816 87012 19820 87068
rect 19820 87012 19876 87068
rect 19876 87012 19880 87068
rect 19816 87008 19880 87012
rect 50296 87068 50360 87072
rect 50296 87012 50300 87068
rect 50300 87012 50356 87068
rect 50356 87012 50360 87068
rect 50296 87008 50360 87012
rect 50376 87068 50440 87072
rect 50376 87012 50380 87068
rect 50380 87012 50436 87068
rect 50436 87012 50440 87068
rect 50376 87008 50440 87012
rect 50456 87068 50520 87072
rect 50456 87012 50460 87068
rect 50460 87012 50516 87068
rect 50516 87012 50520 87068
rect 50456 87008 50520 87012
rect 50536 87068 50600 87072
rect 50536 87012 50540 87068
rect 50540 87012 50596 87068
rect 50596 87012 50600 87068
rect 50536 87008 50600 87012
rect 4216 86524 4280 86528
rect 4216 86468 4220 86524
rect 4220 86468 4276 86524
rect 4276 86468 4280 86524
rect 4216 86464 4280 86468
rect 4296 86524 4360 86528
rect 4296 86468 4300 86524
rect 4300 86468 4356 86524
rect 4356 86468 4360 86524
rect 4296 86464 4360 86468
rect 4376 86524 4440 86528
rect 4376 86468 4380 86524
rect 4380 86468 4436 86524
rect 4436 86468 4440 86524
rect 4376 86464 4440 86468
rect 4456 86524 4520 86528
rect 4456 86468 4460 86524
rect 4460 86468 4516 86524
rect 4516 86468 4520 86524
rect 4456 86464 4520 86468
rect 34936 86524 35000 86528
rect 34936 86468 34940 86524
rect 34940 86468 34996 86524
rect 34996 86468 35000 86524
rect 34936 86464 35000 86468
rect 35016 86524 35080 86528
rect 35016 86468 35020 86524
rect 35020 86468 35076 86524
rect 35076 86468 35080 86524
rect 35016 86464 35080 86468
rect 35096 86524 35160 86528
rect 35096 86468 35100 86524
rect 35100 86468 35156 86524
rect 35156 86468 35160 86524
rect 35096 86464 35160 86468
rect 35176 86524 35240 86528
rect 35176 86468 35180 86524
rect 35180 86468 35236 86524
rect 35236 86468 35240 86524
rect 35176 86464 35240 86468
rect 65656 86524 65720 86528
rect 65656 86468 65660 86524
rect 65660 86468 65716 86524
rect 65716 86468 65720 86524
rect 65656 86464 65720 86468
rect 65736 86524 65800 86528
rect 65736 86468 65740 86524
rect 65740 86468 65796 86524
rect 65796 86468 65800 86524
rect 65736 86464 65800 86468
rect 65816 86524 65880 86528
rect 65816 86468 65820 86524
rect 65820 86468 65876 86524
rect 65876 86468 65880 86524
rect 65816 86464 65880 86468
rect 65896 86524 65960 86528
rect 65896 86468 65900 86524
rect 65900 86468 65956 86524
rect 65956 86468 65960 86524
rect 65896 86464 65960 86468
rect 19576 85980 19640 85984
rect 19576 85924 19580 85980
rect 19580 85924 19636 85980
rect 19636 85924 19640 85980
rect 19576 85920 19640 85924
rect 19656 85980 19720 85984
rect 19656 85924 19660 85980
rect 19660 85924 19716 85980
rect 19716 85924 19720 85980
rect 19656 85920 19720 85924
rect 19736 85980 19800 85984
rect 19736 85924 19740 85980
rect 19740 85924 19796 85980
rect 19796 85924 19800 85980
rect 19736 85920 19800 85924
rect 19816 85980 19880 85984
rect 19816 85924 19820 85980
rect 19820 85924 19876 85980
rect 19876 85924 19880 85980
rect 19816 85920 19880 85924
rect 50296 85980 50360 85984
rect 50296 85924 50300 85980
rect 50300 85924 50356 85980
rect 50356 85924 50360 85980
rect 50296 85920 50360 85924
rect 50376 85980 50440 85984
rect 50376 85924 50380 85980
rect 50380 85924 50436 85980
rect 50436 85924 50440 85980
rect 50376 85920 50440 85924
rect 50456 85980 50520 85984
rect 50456 85924 50460 85980
rect 50460 85924 50516 85980
rect 50516 85924 50520 85980
rect 50456 85920 50520 85924
rect 50536 85980 50600 85984
rect 50536 85924 50540 85980
rect 50540 85924 50596 85980
rect 50596 85924 50600 85980
rect 50536 85920 50600 85924
rect 4216 85436 4280 85440
rect 4216 85380 4220 85436
rect 4220 85380 4276 85436
rect 4276 85380 4280 85436
rect 4216 85376 4280 85380
rect 4296 85436 4360 85440
rect 4296 85380 4300 85436
rect 4300 85380 4356 85436
rect 4356 85380 4360 85436
rect 4296 85376 4360 85380
rect 4376 85436 4440 85440
rect 4376 85380 4380 85436
rect 4380 85380 4436 85436
rect 4436 85380 4440 85436
rect 4376 85376 4440 85380
rect 4456 85436 4520 85440
rect 4456 85380 4460 85436
rect 4460 85380 4516 85436
rect 4516 85380 4520 85436
rect 4456 85376 4520 85380
rect 34936 85436 35000 85440
rect 34936 85380 34940 85436
rect 34940 85380 34996 85436
rect 34996 85380 35000 85436
rect 34936 85376 35000 85380
rect 35016 85436 35080 85440
rect 35016 85380 35020 85436
rect 35020 85380 35076 85436
rect 35076 85380 35080 85436
rect 35016 85376 35080 85380
rect 35096 85436 35160 85440
rect 35096 85380 35100 85436
rect 35100 85380 35156 85436
rect 35156 85380 35160 85436
rect 35096 85376 35160 85380
rect 35176 85436 35240 85440
rect 35176 85380 35180 85436
rect 35180 85380 35236 85436
rect 35236 85380 35240 85436
rect 35176 85376 35240 85380
rect 65656 85436 65720 85440
rect 65656 85380 65660 85436
rect 65660 85380 65716 85436
rect 65716 85380 65720 85436
rect 65656 85376 65720 85380
rect 65736 85436 65800 85440
rect 65736 85380 65740 85436
rect 65740 85380 65796 85436
rect 65796 85380 65800 85436
rect 65736 85376 65800 85380
rect 65816 85436 65880 85440
rect 65816 85380 65820 85436
rect 65820 85380 65876 85436
rect 65876 85380 65880 85436
rect 65816 85376 65880 85380
rect 65896 85436 65960 85440
rect 65896 85380 65900 85436
rect 65900 85380 65956 85436
rect 65956 85380 65960 85436
rect 65896 85376 65960 85380
rect 19576 84892 19640 84896
rect 19576 84836 19580 84892
rect 19580 84836 19636 84892
rect 19636 84836 19640 84892
rect 19576 84832 19640 84836
rect 19656 84892 19720 84896
rect 19656 84836 19660 84892
rect 19660 84836 19716 84892
rect 19716 84836 19720 84892
rect 19656 84832 19720 84836
rect 19736 84892 19800 84896
rect 19736 84836 19740 84892
rect 19740 84836 19796 84892
rect 19796 84836 19800 84892
rect 19736 84832 19800 84836
rect 19816 84892 19880 84896
rect 19816 84836 19820 84892
rect 19820 84836 19876 84892
rect 19876 84836 19880 84892
rect 19816 84832 19880 84836
rect 50296 84892 50360 84896
rect 50296 84836 50300 84892
rect 50300 84836 50356 84892
rect 50356 84836 50360 84892
rect 50296 84832 50360 84836
rect 50376 84892 50440 84896
rect 50376 84836 50380 84892
rect 50380 84836 50436 84892
rect 50436 84836 50440 84892
rect 50376 84832 50440 84836
rect 50456 84892 50520 84896
rect 50456 84836 50460 84892
rect 50460 84836 50516 84892
rect 50516 84836 50520 84892
rect 50456 84832 50520 84836
rect 50536 84892 50600 84896
rect 50536 84836 50540 84892
rect 50540 84836 50596 84892
rect 50596 84836 50600 84892
rect 50536 84832 50600 84836
rect 4216 84348 4280 84352
rect 4216 84292 4220 84348
rect 4220 84292 4276 84348
rect 4276 84292 4280 84348
rect 4216 84288 4280 84292
rect 4296 84348 4360 84352
rect 4296 84292 4300 84348
rect 4300 84292 4356 84348
rect 4356 84292 4360 84348
rect 4296 84288 4360 84292
rect 4376 84348 4440 84352
rect 4376 84292 4380 84348
rect 4380 84292 4436 84348
rect 4436 84292 4440 84348
rect 4376 84288 4440 84292
rect 4456 84348 4520 84352
rect 4456 84292 4460 84348
rect 4460 84292 4516 84348
rect 4516 84292 4520 84348
rect 4456 84288 4520 84292
rect 34936 84348 35000 84352
rect 34936 84292 34940 84348
rect 34940 84292 34996 84348
rect 34996 84292 35000 84348
rect 34936 84288 35000 84292
rect 35016 84348 35080 84352
rect 35016 84292 35020 84348
rect 35020 84292 35076 84348
rect 35076 84292 35080 84348
rect 35016 84288 35080 84292
rect 35096 84348 35160 84352
rect 35096 84292 35100 84348
rect 35100 84292 35156 84348
rect 35156 84292 35160 84348
rect 35096 84288 35160 84292
rect 35176 84348 35240 84352
rect 35176 84292 35180 84348
rect 35180 84292 35236 84348
rect 35236 84292 35240 84348
rect 35176 84288 35240 84292
rect 65656 84348 65720 84352
rect 65656 84292 65660 84348
rect 65660 84292 65716 84348
rect 65716 84292 65720 84348
rect 65656 84288 65720 84292
rect 65736 84348 65800 84352
rect 65736 84292 65740 84348
rect 65740 84292 65796 84348
rect 65796 84292 65800 84348
rect 65736 84288 65800 84292
rect 65816 84348 65880 84352
rect 65816 84292 65820 84348
rect 65820 84292 65876 84348
rect 65876 84292 65880 84348
rect 65816 84288 65880 84292
rect 65896 84348 65960 84352
rect 65896 84292 65900 84348
rect 65900 84292 65956 84348
rect 65956 84292 65960 84348
rect 65896 84288 65960 84292
rect 19576 83804 19640 83808
rect 19576 83748 19580 83804
rect 19580 83748 19636 83804
rect 19636 83748 19640 83804
rect 19576 83744 19640 83748
rect 19656 83804 19720 83808
rect 19656 83748 19660 83804
rect 19660 83748 19716 83804
rect 19716 83748 19720 83804
rect 19656 83744 19720 83748
rect 19736 83804 19800 83808
rect 19736 83748 19740 83804
rect 19740 83748 19796 83804
rect 19796 83748 19800 83804
rect 19736 83744 19800 83748
rect 19816 83804 19880 83808
rect 19816 83748 19820 83804
rect 19820 83748 19876 83804
rect 19876 83748 19880 83804
rect 19816 83744 19880 83748
rect 50296 83804 50360 83808
rect 50296 83748 50300 83804
rect 50300 83748 50356 83804
rect 50356 83748 50360 83804
rect 50296 83744 50360 83748
rect 50376 83804 50440 83808
rect 50376 83748 50380 83804
rect 50380 83748 50436 83804
rect 50436 83748 50440 83804
rect 50376 83744 50440 83748
rect 50456 83804 50520 83808
rect 50456 83748 50460 83804
rect 50460 83748 50516 83804
rect 50516 83748 50520 83804
rect 50456 83744 50520 83748
rect 50536 83804 50600 83808
rect 50536 83748 50540 83804
rect 50540 83748 50596 83804
rect 50596 83748 50600 83804
rect 50536 83744 50600 83748
rect 4216 83260 4280 83264
rect 4216 83204 4220 83260
rect 4220 83204 4276 83260
rect 4276 83204 4280 83260
rect 4216 83200 4280 83204
rect 4296 83260 4360 83264
rect 4296 83204 4300 83260
rect 4300 83204 4356 83260
rect 4356 83204 4360 83260
rect 4296 83200 4360 83204
rect 4376 83260 4440 83264
rect 4376 83204 4380 83260
rect 4380 83204 4436 83260
rect 4436 83204 4440 83260
rect 4376 83200 4440 83204
rect 4456 83260 4520 83264
rect 4456 83204 4460 83260
rect 4460 83204 4516 83260
rect 4516 83204 4520 83260
rect 4456 83200 4520 83204
rect 34936 83260 35000 83264
rect 34936 83204 34940 83260
rect 34940 83204 34996 83260
rect 34996 83204 35000 83260
rect 34936 83200 35000 83204
rect 35016 83260 35080 83264
rect 35016 83204 35020 83260
rect 35020 83204 35076 83260
rect 35076 83204 35080 83260
rect 35016 83200 35080 83204
rect 35096 83260 35160 83264
rect 35096 83204 35100 83260
rect 35100 83204 35156 83260
rect 35156 83204 35160 83260
rect 35096 83200 35160 83204
rect 35176 83260 35240 83264
rect 35176 83204 35180 83260
rect 35180 83204 35236 83260
rect 35236 83204 35240 83260
rect 35176 83200 35240 83204
rect 65656 83260 65720 83264
rect 65656 83204 65660 83260
rect 65660 83204 65716 83260
rect 65716 83204 65720 83260
rect 65656 83200 65720 83204
rect 65736 83260 65800 83264
rect 65736 83204 65740 83260
rect 65740 83204 65796 83260
rect 65796 83204 65800 83260
rect 65736 83200 65800 83204
rect 65816 83260 65880 83264
rect 65816 83204 65820 83260
rect 65820 83204 65876 83260
rect 65876 83204 65880 83260
rect 65816 83200 65880 83204
rect 65896 83260 65960 83264
rect 65896 83204 65900 83260
rect 65900 83204 65956 83260
rect 65956 83204 65960 83260
rect 65896 83200 65960 83204
rect 19576 82716 19640 82720
rect 19576 82660 19580 82716
rect 19580 82660 19636 82716
rect 19636 82660 19640 82716
rect 19576 82656 19640 82660
rect 19656 82716 19720 82720
rect 19656 82660 19660 82716
rect 19660 82660 19716 82716
rect 19716 82660 19720 82716
rect 19656 82656 19720 82660
rect 19736 82716 19800 82720
rect 19736 82660 19740 82716
rect 19740 82660 19796 82716
rect 19796 82660 19800 82716
rect 19736 82656 19800 82660
rect 19816 82716 19880 82720
rect 19816 82660 19820 82716
rect 19820 82660 19876 82716
rect 19876 82660 19880 82716
rect 19816 82656 19880 82660
rect 50296 82716 50360 82720
rect 50296 82660 50300 82716
rect 50300 82660 50356 82716
rect 50356 82660 50360 82716
rect 50296 82656 50360 82660
rect 50376 82716 50440 82720
rect 50376 82660 50380 82716
rect 50380 82660 50436 82716
rect 50436 82660 50440 82716
rect 50376 82656 50440 82660
rect 50456 82716 50520 82720
rect 50456 82660 50460 82716
rect 50460 82660 50516 82716
rect 50516 82660 50520 82716
rect 50456 82656 50520 82660
rect 50536 82716 50600 82720
rect 50536 82660 50540 82716
rect 50540 82660 50596 82716
rect 50596 82660 50600 82716
rect 50536 82656 50600 82660
rect 4216 82172 4280 82176
rect 4216 82116 4220 82172
rect 4220 82116 4276 82172
rect 4276 82116 4280 82172
rect 4216 82112 4280 82116
rect 4296 82172 4360 82176
rect 4296 82116 4300 82172
rect 4300 82116 4356 82172
rect 4356 82116 4360 82172
rect 4296 82112 4360 82116
rect 4376 82172 4440 82176
rect 4376 82116 4380 82172
rect 4380 82116 4436 82172
rect 4436 82116 4440 82172
rect 4376 82112 4440 82116
rect 4456 82172 4520 82176
rect 4456 82116 4460 82172
rect 4460 82116 4516 82172
rect 4516 82116 4520 82172
rect 4456 82112 4520 82116
rect 34936 82172 35000 82176
rect 34936 82116 34940 82172
rect 34940 82116 34996 82172
rect 34996 82116 35000 82172
rect 34936 82112 35000 82116
rect 35016 82172 35080 82176
rect 35016 82116 35020 82172
rect 35020 82116 35076 82172
rect 35076 82116 35080 82172
rect 35016 82112 35080 82116
rect 35096 82172 35160 82176
rect 35096 82116 35100 82172
rect 35100 82116 35156 82172
rect 35156 82116 35160 82172
rect 35096 82112 35160 82116
rect 35176 82172 35240 82176
rect 35176 82116 35180 82172
rect 35180 82116 35236 82172
rect 35236 82116 35240 82172
rect 35176 82112 35240 82116
rect 65656 82172 65720 82176
rect 65656 82116 65660 82172
rect 65660 82116 65716 82172
rect 65716 82116 65720 82172
rect 65656 82112 65720 82116
rect 65736 82172 65800 82176
rect 65736 82116 65740 82172
rect 65740 82116 65796 82172
rect 65796 82116 65800 82172
rect 65736 82112 65800 82116
rect 65816 82172 65880 82176
rect 65816 82116 65820 82172
rect 65820 82116 65876 82172
rect 65876 82116 65880 82172
rect 65816 82112 65880 82116
rect 65896 82172 65960 82176
rect 65896 82116 65900 82172
rect 65900 82116 65956 82172
rect 65956 82116 65960 82172
rect 65896 82112 65960 82116
rect 19576 81628 19640 81632
rect 19576 81572 19580 81628
rect 19580 81572 19636 81628
rect 19636 81572 19640 81628
rect 19576 81568 19640 81572
rect 19656 81628 19720 81632
rect 19656 81572 19660 81628
rect 19660 81572 19716 81628
rect 19716 81572 19720 81628
rect 19656 81568 19720 81572
rect 19736 81628 19800 81632
rect 19736 81572 19740 81628
rect 19740 81572 19796 81628
rect 19796 81572 19800 81628
rect 19736 81568 19800 81572
rect 19816 81628 19880 81632
rect 19816 81572 19820 81628
rect 19820 81572 19876 81628
rect 19876 81572 19880 81628
rect 19816 81568 19880 81572
rect 50296 81628 50360 81632
rect 50296 81572 50300 81628
rect 50300 81572 50356 81628
rect 50356 81572 50360 81628
rect 50296 81568 50360 81572
rect 50376 81628 50440 81632
rect 50376 81572 50380 81628
rect 50380 81572 50436 81628
rect 50436 81572 50440 81628
rect 50376 81568 50440 81572
rect 50456 81628 50520 81632
rect 50456 81572 50460 81628
rect 50460 81572 50516 81628
rect 50516 81572 50520 81628
rect 50456 81568 50520 81572
rect 50536 81628 50600 81632
rect 50536 81572 50540 81628
rect 50540 81572 50596 81628
rect 50596 81572 50600 81628
rect 50536 81568 50600 81572
rect 4216 81084 4280 81088
rect 4216 81028 4220 81084
rect 4220 81028 4276 81084
rect 4276 81028 4280 81084
rect 4216 81024 4280 81028
rect 4296 81084 4360 81088
rect 4296 81028 4300 81084
rect 4300 81028 4356 81084
rect 4356 81028 4360 81084
rect 4296 81024 4360 81028
rect 4376 81084 4440 81088
rect 4376 81028 4380 81084
rect 4380 81028 4436 81084
rect 4436 81028 4440 81084
rect 4376 81024 4440 81028
rect 4456 81084 4520 81088
rect 4456 81028 4460 81084
rect 4460 81028 4516 81084
rect 4516 81028 4520 81084
rect 4456 81024 4520 81028
rect 34936 81084 35000 81088
rect 34936 81028 34940 81084
rect 34940 81028 34996 81084
rect 34996 81028 35000 81084
rect 34936 81024 35000 81028
rect 35016 81084 35080 81088
rect 35016 81028 35020 81084
rect 35020 81028 35076 81084
rect 35076 81028 35080 81084
rect 35016 81024 35080 81028
rect 35096 81084 35160 81088
rect 35096 81028 35100 81084
rect 35100 81028 35156 81084
rect 35156 81028 35160 81084
rect 35096 81024 35160 81028
rect 35176 81084 35240 81088
rect 35176 81028 35180 81084
rect 35180 81028 35236 81084
rect 35236 81028 35240 81084
rect 35176 81024 35240 81028
rect 65656 81084 65720 81088
rect 65656 81028 65660 81084
rect 65660 81028 65716 81084
rect 65716 81028 65720 81084
rect 65656 81024 65720 81028
rect 65736 81084 65800 81088
rect 65736 81028 65740 81084
rect 65740 81028 65796 81084
rect 65796 81028 65800 81084
rect 65736 81024 65800 81028
rect 65816 81084 65880 81088
rect 65816 81028 65820 81084
rect 65820 81028 65876 81084
rect 65876 81028 65880 81084
rect 65816 81024 65880 81028
rect 65896 81084 65960 81088
rect 65896 81028 65900 81084
rect 65900 81028 65956 81084
rect 65956 81028 65960 81084
rect 65896 81024 65960 81028
rect 19576 80540 19640 80544
rect 19576 80484 19580 80540
rect 19580 80484 19636 80540
rect 19636 80484 19640 80540
rect 19576 80480 19640 80484
rect 19656 80540 19720 80544
rect 19656 80484 19660 80540
rect 19660 80484 19716 80540
rect 19716 80484 19720 80540
rect 19656 80480 19720 80484
rect 19736 80540 19800 80544
rect 19736 80484 19740 80540
rect 19740 80484 19796 80540
rect 19796 80484 19800 80540
rect 19736 80480 19800 80484
rect 19816 80540 19880 80544
rect 19816 80484 19820 80540
rect 19820 80484 19876 80540
rect 19876 80484 19880 80540
rect 19816 80480 19880 80484
rect 50296 80540 50360 80544
rect 50296 80484 50300 80540
rect 50300 80484 50356 80540
rect 50356 80484 50360 80540
rect 50296 80480 50360 80484
rect 50376 80540 50440 80544
rect 50376 80484 50380 80540
rect 50380 80484 50436 80540
rect 50436 80484 50440 80540
rect 50376 80480 50440 80484
rect 50456 80540 50520 80544
rect 50456 80484 50460 80540
rect 50460 80484 50516 80540
rect 50516 80484 50520 80540
rect 50456 80480 50520 80484
rect 50536 80540 50600 80544
rect 50536 80484 50540 80540
rect 50540 80484 50596 80540
rect 50596 80484 50600 80540
rect 50536 80480 50600 80484
rect 4216 79996 4280 80000
rect 4216 79940 4220 79996
rect 4220 79940 4276 79996
rect 4276 79940 4280 79996
rect 4216 79936 4280 79940
rect 4296 79996 4360 80000
rect 4296 79940 4300 79996
rect 4300 79940 4356 79996
rect 4356 79940 4360 79996
rect 4296 79936 4360 79940
rect 4376 79996 4440 80000
rect 4376 79940 4380 79996
rect 4380 79940 4436 79996
rect 4436 79940 4440 79996
rect 4376 79936 4440 79940
rect 4456 79996 4520 80000
rect 4456 79940 4460 79996
rect 4460 79940 4516 79996
rect 4516 79940 4520 79996
rect 4456 79936 4520 79940
rect 34936 79996 35000 80000
rect 34936 79940 34940 79996
rect 34940 79940 34996 79996
rect 34996 79940 35000 79996
rect 34936 79936 35000 79940
rect 35016 79996 35080 80000
rect 35016 79940 35020 79996
rect 35020 79940 35076 79996
rect 35076 79940 35080 79996
rect 35016 79936 35080 79940
rect 35096 79996 35160 80000
rect 35096 79940 35100 79996
rect 35100 79940 35156 79996
rect 35156 79940 35160 79996
rect 35096 79936 35160 79940
rect 35176 79996 35240 80000
rect 35176 79940 35180 79996
rect 35180 79940 35236 79996
rect 35236 79940 35240 79996
rect 35176 79936 35240 79940
rect 65656 79996 65720 80000
rect 65656 79940 65660 79996
rect 65660 79940 65716 79996
rect 65716 79940 65720 79996
rect 65656 79936 65720 79940
rect 65736 79996 65800 80000
rect 65736 79940 65740 79996
rect 65740 79940 65796 79996
rect 65796 79940 65800 79996
rect 65736 79936 65800 79940
rect 65816 79996 65880 80000
rect 65816 79940 65820 79996
rect 65820 79940 65876 79996
rect 65876 79940 65880 79996
rect 65816 79936 65880 79940
rect 65896 79996 65960 80000
rect 65896 79940 65900 79996
rect 65900 79940 65956 79996
rect 65956 79940 65960 79996
rect 65896 79936 65960 79940
rect 19576 79452 19640 79456
rect 19576 79396 19580 79452
rect 19580 79396 19636 79452
rect 19636 79396 19640 79452
rect 19576 79392 19640 79396
rect 19656 79452 19720 79456
rect 19656 79396 19660 79452
rect 19660 79396 19716 79452
rect 19716 79396 19720 79452
rect 19656 79392 19720 79396
rect 19736 79452 19800 79456
rect 19736 79396 19740 79452
rect 19740 79396 19796 79452
rect 19796 79396 19800 79452
rect 19736 79392 19800 79396
rect 19816 79452 19880 79456
rect 19816 79396 19820 79452
rect 19820 79396 19876 79452
rect 19876 79396 19880 79452
rect 19816 79392 19880 79396
rect 50296 79452 50360 79456
rect 50296 79396 50300 79452
rect 50300 79396 50356 79452
rect 50356 79396 50360 79452
rect 50296 79392 50360 79396
rect 50376 79452 50440 79456
rect 50376 79396 50380 79452
rect 50380 79396 50436 79452
rect 50436 79396 50440 79452
rect 50376 79392 50440 79396
rect 50456 79452 50520 79456
rect 50456 79396 50460 79452
rect 50460 79396 50516 79452
rect 50516 79396 50520 79452
rect 50456 79392 50520 79396
rect 50536 79452 50600 79456
rect 50536 79396 50540 79452
rect 50540 79396 50596 79452
rect 50596 79396 50600 79452
rect 50536 79392 50600 79396
rect 4216 78908 4280 78912
rect 4216 78852 4220 78908
rect 4220 78852 4276 78908
rect 4276 78852 4280 78908
rect 4216 78848 4280 78852
rect 4296 78908 4360 78912
rect 4296 78852 4300 78908
rect 4300 78852 4356 78908
rect 4356 78852 4360 78908
rect 4296 78848 4360 78852
rect 4376 78908 4440 78912
rect 4376 78852 4380 78908
rect 4380 78852 4436 78908
rect 4436 78852 4440 78908
rect 4376 78848 4440 78852
rect 4456 78908 4520 78912
rect 4456 78852 4460 78908
rect 4460 78852 4516 78908
rect 4516 78852 4520 78908
rect 4456 78848 4520 78852
rect 34936 78908 35000 78912
rect 34936 78852 34940 78908
rect 34940 78852 34996 78908
rect 34996 78852 35000 78908
rect 34936 78848 35000 78852
rect 35016 78908 35080 78912
rect 35016 78852 35020 78908
rect 35020 78852 35076 78908
rect 35076 78852 35080 78908
rect 35016 78848 35080 78852
rect 35096 78908 35160 78912
rect 35096 78852 35100 78908
rect 35100 78852 35156 78908
rect 35156 78852 35160 78908
rect 35096 78848 35160 78852
rect 35176 78908 35240 78912
rect 35176 78852 35180 78908
rect 35180 78852 35236 78908
rect 35236 78852 35240 78908
rect 35176 78848 35240 78852
rect 65656 78908 65720 78912
rect 65656 78852 65660 78908
rect 65660 78852 65716 78908
rect 65716 78852 65720 78908
rect 65656 78848 65720 78852
rect 65736 78908 65800 78912
rect 65736 78852 65740 78908
rect 65740 78852 65796 78908
rect 65796 78852 65800 78908
rect 65736 78848 65800 78852
rect 65816 78908 65880 78912
rect 65816 78852 65820 78908
rect 65820 78852 65876 78908
rect 65876 78852 65880 78908
rect 65816 78848 65880 78852
rect 65896 78908 65960 78912
rect 65896 78852 65900 78908
rect 65900 78852 65956 78908
rect 65956 78852 65960 78908
rect 65896 78848 65960 78852
rect 19576 78364 19640 78368
rect 19576 78308 19580 78364
rect 19580 78308 19636 78364
rect 19636 78308 19640 78364
rect 19576 78304 19640 78308
rect 19656 78364 19720 78368
rect 19656 78308 19660 78364
rect 19660 78308 19716 78364
rect 19716 78308 19720 78364
rect 19656 78304 19720 78308
rect 19736 78364 19800 78368
rect 19736 78308 19740 78364
rect 19740 78308 19796 78364
rect 19796 78308 19800 78364
rect 19736 78304 19800 78308
rect 19816 78364 19880 78368
rect 19816 78308 19820 78364
rect 19820 78308 19876 78364
rect 19876 78308 19880 78364
rect 19816 78304 19880 78308
rect 50296 78364 50360 78368
rect 50296 78308 50300 78364
rect 50300 78308 50356 78364
rect 50356 78308 50360 78364
rect 50296 78304 50360 78308
rect 50376 78364 50440 78368
rect 50376 78308 50380 78364
rect 50380 78308 50436 78364
rect 50436 78308 50440 78364
rect 50376 78304 50440 78308
rect 50456 78364 50520 78368
rect 50456 78308 50460 78364
rect 50460 78308 50516 78364
rect 50516 78308 50520 78364
rect 50456 78304 50520 78308
rect 50536 78364 50600 78368
rect 50536 78308 50540 78364
rect 50540 78308 50596 78364
rect 50596 78308 50600 78364
rect 50536 78304 50600 78308
rect 4216 77820 4280 77824
rect 4216 77764 4220 77820
rect 4220 77764 4276 77820
rect 4276 77764 4280 77820
rect 4216 77760 4280 77764
rect 4296 77820 4360 77824
rect 4296 77764 4300 77820
rect 4300 77764 4356 77820
rect 4356 77764 4360 77820
rect 4296 77760 4360 77764
rect 4376 77820 4440 77824
rect 4376 77764 4380 77820
rect 4380 77764 4436 77820
rect 4436 77764 4440 77820
rect 4376 77760 4440 77764
rect 4456 77820 4520 77824
rect 4456 77764 4460 77820
rect 4460 77764 4516 77820
rect 4516 77764 4520 77820
rect 4456 77760 4520 77764
rect 34936 77820 35000 77824
rect 34936 77764 34940 77820
rect 34940 77764 34996 77820
rect 34996 77764 35000 77820
rect 34936 77760 35000 77764
rect 35016 77820 35080 77824
rect 35016 77764 35020 77820
rect 35020 77764 35076 77820
rect 35076 77764 35080 77820
rect 35016 77760 35080 77764
rect 35096 77820 35160 77824
rect 35096 77764 35100 77820
rect 35100 77764 35156 77820
rect 35156 77764 35160 77820
rect 35096 77760 35160 77764
rect 35176 77820 35240 77824
rect 35176 77764 35180 77820
rect 35180 77764 35236 77820
rect 35236 77764 35240 77820
rect 35176 77760 35240 77764
rect 65656 77820 65720 77824
rect 65656 77764 65660 77820
rect 65660 77764 65716 77820
rect 65716 77764 65720 77820
rect 65656 77760 65720 77764
rect 65736 77820 65800 77824
rect 65736 77764 65740 77820
rect 65740 77764 65796 77820
rect 65796 77764 65800 77820
rect 65736 77760 65800 77764
rect 65816 77820 65880 77824
rect 65816 77764 65820 77820
rect 65820 77764 65876 77820
rect 65876 77764 65880 77820
rect 65816 77760 65880 77764
rect 65896 77820 65960 77824
rect 65896 77764 65900 77820
rect 65900 77764 65956 77820
rect 65956 77764 65960 77820
rect 65896 77760 65960 77764
rect 19576 77276 19640 77280
rect 19576 77220 19580 77276
rect 19580 77220 19636 77276
rect 19636 77220 19640 77276
rect 19576 77216 19640 77220
rect 19656 77276 19720 77280
rect 19656 77220 19660 77276
rect 19660 77220 19716 77276
rect 19716 77220 19720 77276
rect 19656 77216 19720 77220
rect 19736 77276 19800 77280
rect 19736 77220 19740 77276
rect 19740 77220 19796 77276
rect 19796 77220 19800 77276
rect 19736 77216 19800 77220
rect 19816 77276 19880 77280
rect 19816 77220 19820 77276
rect 19820 77220 19876 77276
rect 19876 77220 19880 77276
rect 19816 77216 19880 77220
rect 50296 77276 50360 77280
rect 50296 77220 50300 77276
rect 50300 77220 50356 77276
rect 50356 77220 50360 77276
rect 50296 77216 50360 77220
rect 50376 77276 50440 77280
rect 50376 77220 50380 77276
rect 50380 77220 50436 77276
rect 50436 77220 50440 77276
rect 50376 77216 50440 77220
rect 50456 77276 50520 77280
rect 50456 77220 50460 77276
rect 50460 77220 50516 77276
rect 50516 77220 50520 77276
rect 50456 77216 50520 77220
rect 50536 77276 50600 77280
rect 50536 77220 50540 77276
rect 50540 77220 50596 77276
rect 50596 77220 50600 77276
rect 50536 77216 50600 77220
rect 4216 76732 4280 76736
rect 4216 76676 4220 76732
rect 4220 76676 4276 76732
rect 4276 76676 4280 76732
rect 4216 76672 4280 76676
rect 4296 76732 4360 76736
rect 4296 76676 4300 76732
rect 4300 76676 4356 76732
rect 4356 76676 4360 76732
rect 4296 76672 4360 76676
rect 4376 76732 4440 76736
rect 4376 76676 4380 76732
rect 4380 76676 4436 76732
rect 4436 76676 4440 76732
rect 4376 76672 4440 76676
rect 4456 76732 4520 76736
rect 4456 76676 4460 76732
rect 4460 76676 4516 76732
rect 4516 76676 4520 76732
rect 4456 76672 4520 76676
rect 34936 76732 35000 76736
rect 34936 76676 34940 76732
rect 34940 76676 34996 76732
rect 34996 76676 35000 76732
rect 34936 76672 35000 76676
rect 35016 76732 35080 76736
rect 35016 76676 35020 76732
rect 35020 76676 35076 76732
rect 35076 76676 35080 76732
rect 35016 76672 35080 76676
rect 35096 76732 35160 76736
rect 35096 76676 35100 76732
rect 35100 76676 35156 76732
rect 35156 76676 35160 76732
rect 35096 76672 35160 76676
rect 35176 76732 35240 76736
rect 35176 76676 35180 76732
rect 35180 76676 35236 76732
rect 35236 76676 35240 76732
rect 35176 76672 35240 76676
rect 65656 76732 65720 76736
rect 65656 76676 65660 76732
rect 65660 76676 65716 76732
rect 65716 76676 65720 76732
rect 65656 76672 65720 76676
rect 65736 76732 65800 76736
rect 65736 76676 65740 76732
rect 65740 76676 65796 76732
rect 65796 76676 65800 76732
rect 65736 76672 65800 76676
rect 65816 76732 65880 76736
rect 65816 76676 65820 76732
rect 65820 76676 65876 76732
rect 65876 76676 65880 76732
rect 65816 76672 65880 76676
rect 65896 76732 65960 76736
rect 65896 76676 65900 76732
rect 65900 76676 65956 76732
rect 65956 76676 65960 76732
rect 65896 76672 65960 76676
rect 19576 76188 19640 76192
rect 19576 76132 19580 76188
rect 19580 76132 19636 76188
rect 19636 76132 19640 76188
rect 19576 76128 19640 76132
rect 19656 76188 19720 76192
rect 19656 76132 19660 76188
rect 19660 76132 19716 76188
rect 19716 76132 19720 76188
rect 19656 76128 19720 76132
rect 19736 76188 19800 76192
rect 19736 76132 19740 76188
rect 19740 76132 19796 76188
rect 19796 76132 19800 76188
rect 19736 76128 19800 76132
rect 19816 76188 19880 76192
rect 19816 76132 19820 76188
rect 19820 76132 19876 76188
rect 19876 76132 19880 76188
rect 19816 76128 19880 76132
rect 50296 76188 50360 76192
rect 50296 76132 50300 76188
rect 50300 76132 50356 76188
rect 50356 76132 50360 76188
rect 50296 76128 50360 76132
rect 50376 76188 50440 76192
rect 50376 76132 50380 76188
rect 50380 76132 50436 76188
rect 50436 76132 50440 76188
rect 50376 76128 50440 76132
rect 50456 76188 50520 76192
rect 50456 76132 50460 76188
rect 50460 76132 50516 76188
rect 50516 76132 50520 76188
rect 50456 76128 50520 76132
rect 50536 76188 50600 76192
rect 50536 76132 50540 76188
rect 50540 76132 50596 76188
rect 50596 76132 50600 76188
rect 50536 76128 50600 76132
rect 4216 75644 4280 75648
rect 4216 75588 4220 75644
rect 4220 75588 4276 75644
rect 4276 75588 4280 75644
rect 4216 75584 4280 75588
rect 4296 75644 4360 75648
rect 4296 75588 4300 75644
rect 4300 75588 4356 75644
rect 4356 75588 4360 75644
rect 4296 75584 4360 75588
rect 4376 75644 4440 75648
rect 4376 75588 4380 75644
rect 4380 75588 4436 75644
rect 4436 75588 4440 75644
rect 4376 75584 4440 75588
rect 4456 75644 4520 75648
rect 4456 75588 4460 75644
rect 4460 75588 4516 75644
rect 4516 75588 4520 75644
rect 4456 75584 4520 75588
rect 34936 75644 35000 75648
rect 34936 75588 34940 75644
rect 34940 75588 34996 75644
rect 34996 75588 35000 75644
rect 34936 75584 35000 75588
rect 35016 75644 35080 75648
rect 35016 75588 35020 75644
rect 35020 75588 35076 75644
rect 35076 75588 35080 75644
rect 35016 75584 35080 75588
rect 35096 75644 35160 75648
rect 35096 75588 35100 75644
rect 35100 75588 35156 75644
rect 35156 75588 35160 75644
rect 35096 75584 35160 75588
rect 35176 75644 35240 75648
rect 35176 75588 35180 75644
rect 35180 75588 35236 75644
rect 35236 75588 35240 75644
rect 35176 75584 35240 75588
rect 65656 75644 65720 75648
rect 65656 75588 65660 75644
rect 65660 75588 65716 75644
rect 65716 75588 65720 75644
rect 65656 75584 65720 75588
rect 65736 75644 65800 75648
rect 65736 75588 65740 75644
rect 65740 75588 65796 75644
rect 65796 75588 65800 75644
rect 65736 75584 65800 75588
rect 65816 75644 65880 75648
rect 65816 75588 65820 75644
rect 65820 75588 65876 75644
rect 65876 75588 65880 75644
rect 65816 75584 65880 75588
rect 65896 75644 65960 75648
rect 65896 75588 65900 75644
rect 65900 75588 65956 75644
rect 65956 75588 65960 75644
rect 65896 75584 65960 75588
rect 19576 75100 19640 75104
rect 19576 75044 19580 75100
rect 19580 75044 19636 75100
rect 19636 75044 19640 75100
rect 19576 75040 19640 75044
rect 19656 75100 19720 75104
rect 19656 75044 19660 75100
rect 19660 75044 19716 75100
rect 19716 75044 19720 75100
rect 19656 75040 19720 75044
rect 19736 75100 19800 75104
rect 19736 75044 19740 75100
rect 19740 75044 19796 75100
rect 19796 75044 19800 75100
rect 19736 75040 19800 75044
rect 19816 75100 19880 75104
rect 19816 75044 19820 75100
rect 19820 75044 19876 75100
rect 19876 75044 19880 75100
rect 19816 75040 19880 75044
rect 50296 75100 50360 75104
rect 50296 75044 50300 75100
rect 50300 75044 50356 75100
rect 50356 75044 50360 75100
rect 50296 75040 50360 75044
rect 50376 75100 50440 75104
rect 50376 75044 50380 75100
rect 50380 75044 50436 75100
rect 50436 75044 50440 75100
rect 50376 75040 50440 75044
rect 50456 75100 50520 75104
rect 50456 75044 50460 75100
rect 50460 75044 50516 75100
rect 50516 75044 50520 75100
rect 50456 75040 50520 75044
rect 50536 75100 50600 75104
rect 50536 75044 50540 75100
rect 50540 75044 50596 75100
rect 50596 75044 50600 75100
rect 50536 75040 50600 75044
rect 4216 74556 4280 74560
rect 4216 74500 4220 74556
rect 4220 74500 4276 74556
rect 4276 74500 4280 74556
rect 4216 74496 4280 74500
rect 4296 74556 4360 74560
rect 4296 74500 4300 74556
rect 4300 74500 4356 74556
rect 4356 74500 4360 74556
rect 4296 74496 4360 74500
rect 4376 74556 4440 74560
rect 4376 74500 4380 74556
rect 4380 74500 4436 74556
rect 4436 74500 4440 74556
rect 4376 74496 4440 74500
rect 4456 74556 4520 74560
rect 4456 74500 4460 74556
rect 4460 74500 4516 74556
rect 4516 74500 4520 74556
rect 4456 74496 4520 74500
rect 34936 74556 35000 74560
rect 34936 74500 34940 74556
rect 34940 74500 34996 74556
rect 34996 74500 35000 74556
rect 34936 74496 35000 74500
rect 35016 74556 35080 74560
rect 35016 74500 35020 74556
rect 35020 74500 35076 74556
rect 35076 74500 35080 74556
rect 35016 74496 35080 74500
rect 35096 74556 35160 74560
rect 35096 74500 35100 74556
rect 35100 74500 35156 74556
rect 35156 74500 35160 74556
rect 35096 74496 35160 74500
rect 35176 74556 35240 74560
rect 35176 74500 35180 74556
rect 35180 74500 35236 74556
rect 35236 74500 35240 74556
rect 35176 74496 35240 74500
rect 65656 74556 65720 74560
rect 65656 74500 65660 74556
rect 65660 74500 65716 74556
rect 65716 74500 65720 74556
rect 65656 74496 65720 74500
rect 65736 74556 65800 74560
rect 65736 74500 65740 74556
rect 65740 74500 65796 74556
rect 65796 74500 65800 74556
rect 65736 74496 65800 74500
rect 65816 74556 65880 74560
rect 65816 74500 65820 74556
rect 65820 74500 65876 74556
rect 65876 74500 65880 74556
rect 65816 74496 65880 74500
rect 65896 74556 65960 74560
rect 65896 74500 65900 74556
rect 65900 74500 65956 74556
rect 65956 74500 65960 74556
rect 65896 74496 65960 74500
rect 19576 74012 19640 74016
rect 19576 73956 19580 74012
rect 19580 73956 19636 74012
rect 19636 73956 19640 74012
rect 19576 73952 19640 73956
rect 19656 74012 19720 74016
rect 19656 73956 19660 74012
rect 19660 73956 19716 74012
rect 19716 73956 19720 74012
rect 19656 73952 19720 73956
rect 19736 74012 19800 74016
rect 19736 73956 19740 74012
rect 19740 73956 19796 74012
rect 19796 73956 19800 74012
rect 19736 73952 19800 73956
rect 19816 74012 19880 74016
rect 19816 73956 19820 74012
rect 19820 73956 19876 74012
rect 19876 73956 19880 74012
rect 19816 73952 19880 73956
rect 50296 74012 50360 74016
rect 50296 73956 50300 74012
rect 50300 73956 50356 74012
rect 50356 73956 50360 74012
rect 50296 73952 50360 73956
rect 50376 74012 50440 74016
rect 50376 73956 50380 74012
rect 50380 73956 50436 74012
rect 50436 73956 50440 74012
rect 50376 73952 50440 73956
rect 50456 74012 50520 74016
rect 50456 73956 50460 74012
rect 50460 73956 50516 74012
rect 50516 73956 50520 74012
rect 50456 73952 50520 73956
rect 50536 74012 50600 74016
rect 50536 73956 50540 74012
rect 50540 73956 50596 74012
rect 50596 73956 50600 74012
rect 50536 73952 50600 73956
rect 4216 73468 4280 73472
rect 4216 73412 4220 73468
rect 4220 73412 4276 73468
rect 4276 73412 4280 73468
rect 4216 73408 4280 73412
rect 4296 73468 4360 73472
rect 4296 73412 4300 73468
rect 4300 73412 4356 73468
rect 4356 73412 4360 73468
rect 4296 73408 4360 73412
rect 4376 73468 4440 73472
rect 4376 73412 4380 73468
rect 4380 73412 4436 73468
rect 4436 73412 4440 73468
rect 4376 73408 4440 73412
rect 4456 73468 4520 73472
rect 4456 73412 4460 73468
rect 4460 73412 4516 73468
rect 4516 73412 4520 73468
rect 4456 73408 4520 73412
rect 34936 73468 35000 73472
rect 34936 73412 34940 73468
rect 34940 73412 34996 73468
rect 34996 73412 35000 73468
rect 34936 73408 35000 73412
rect 35016 73468 35080 73472
rect 35016 73412 35020 73468
rect 35020 73412 35076 73468
rect 35076 73412 35080 73468
rect 35016 73408 35080 73412
rect 35096 73468 35160 73472
rect 35096 73412 35100 73468
rect 35100 73412 35156 73468
rect 35156 73412 35160 73468
rect 35096 73408 35160 73412
rect 35176 73468 35240 73472
rect 35176 73412 35180 73468
rect 35180 73412 35236 73468
rect 35236 73412 35240 73468
rect 35176 73408 35240 73412
rect 65656 73468 65720 73472
rect 65656 73412 65660 73468
rect 65660 73412 65716 73468
rect 65716 73412 65720 73468
rect 65656 73408 65720 73412
rect 65736 73468 65800 73472
rect 65736 73412 65740 73468
rect 65740 73412 65796 73468
rect 65796 73412 65800 73468
rect 65736 73408 65800 73412
rect 65816 73468 65880 73472
rect 65816 73412 65820 73468
rect 65820 73412 65876 73468
rect 65876 73412 65880 73468
rect 65816 73408 65880 73412
rect 65896 73468 65960 73472
rect 65896 73412 65900 73468
rect 65900 73412 65956 73468
rect 65956 73412 65960 73468
rect 65896 73408 65960 73412
rect 19576 72924 19640 72928
rect 19576 72868 19580 72924
rect 19580 72868 19636 72924
rect 19636 72868 19640 72924
rect 19576 72864 19640 72868
rect 19656 72924 19720 72928
rect 19656 72868 19660 72924
rect 19660 72868 19716 72924
rect 19716 72868 19720 72924
rect 19656 72864 19720 72868
rect 19736 72924 19800 72928
rect 19736 72868 19740 72924
rect 19740 72868 19796 72924
rect 19796 72868 19800 72924
rect 19736 72864 19800 72868
rect 19816 72924 19880 72928
rect 19816 72868 19820 72924
rect 19820 72868 19876 72924
rect 19876 72868 19880 72924
rect 19816 72864 19880 72868
rect 50296 72924 50360 72928
rect 50296 72868 50300 72924
rect 50300 72868 50356 72924
rect 50356 72868 50360 72924
rect 50296 72864 50360 72868
rect 50376 72924 50440 72928
rect 50376 72868 50380 72924
rect 50380 72868 50436 72924
rect 50436 72868 50440 72924
rect 50376 72864 50440 72868
rect 50456 72924 50520 72928
rect 50456 72868 50460 72924
rect 50460 72868 50516 72924
rect 50516 72868 50520 72924
rect 50456 72864 50520 72868
rect 50536 72924 50600 72928
rect 50536 72868 50540 72924
rect 50540 72868 50596 72924
rect 50596 72868 50600 72924
rect 50536 72864 50600 72868
rect 4216 72380 4280 72384
rect 4216 72324 4220 72380
rect 4220 72324 4276 72380
rect 4276 72324 4280 72380
rect 4216 72320 4280 72324
rect 4296 72380 4360 72384
rect 4296 72324 4300 72380
rect 4300 72324 4356 72380
rect 4356 72324 4360 72380
rect 4296 72320 4360 72324
rect 4376 72380 4440 72384
rect 4376 72324 4380 72380
rect 4380 72324 4436 72380
rect 4436 72324 4440 72380
rect 4376 72320 4440 72324
rect 4456 72380 4520 72384
rect 4456 72324 4460 72380
rect 4460 72324 4516 72380
rect 4516 72324 4520 72380
rect 4456 72320 4520 72324
rect 34936 72380 35000 72384
rect 34936 72324 34940 72380
rect 34940 72324 34996 72380
rect 34996 72324 35000 72380
rect 34936 72320 35000 72324
rect 35016 72380 35080 72384
rect 35016 72324 35020 72380
rect 35020 72324 35076 72380
rect 35076 72324 35080 72380
rect 35016 72320 35080 72324
rect 35096 72380 35160 72384
rect 35096 72324 35100 72380
rect 35100 72324 35156 72380
rect 35156 72324 35160 72380
rect 35096 72320 35160 72324
rect 35176 72380 35240 72384
rect 35176 72324 35180 72380
rect 35180 72324 35236 72380
rect 35236 72324 35240 72380
rect 35176 72320 35240 72324
rect 65656 72380 65720 72384
rect 65656 72324 65660 72380
rect 65660 72324 65716 72380
rect 65716 72324 65720 72380
rect 65656 72320 65720 72324
rect 65736 72380 65800 72384
rect 65736 72324 65740 72380
rect 65740 72324 65796 72380
rect 65796 72324 65800 72380
rect 65736 72320 65800 72324
rect 65816 72380 65880 72384
rect 65816 72324 65820 72380
rect 65820 72324 65876 72380
rect 65876 72324 65880 72380
rect 65816 72320 65880 72324
rect 65896 72380 65960 72384
rect 65896 72324 65900 72380
rect 65900 72324 65956 72380
rect 65956 72324 65960 72380
rect 65896 72320 65960 72324
rect 19576 71836 19640 71840
rect 19576 71780 19580 71836
rect 19580 71780 19636 71836
rect 19636 71780 19640 71836
rect 19576 71776 19640 71780
rect 19656 71836 19720 71840
rect 19656 71780 19660 71836
rect 19660 71780 19716 71836
rect 19716 71780 19720 71836
rect 19656 71776 19720 71780
rect 19736 71836 19800 71840
rect 19736 71780 19740 71836
rect 19740 71780 19796 71836
rect 19796 71780 19800 71836
rect 19736 71776 19800 71780
rect 19816 71836 19880 71840
rect 19816 71780 19820 71836
rect 19820 71780 19876 71836
rect 19876 71780 19880 71836
rect 19816 71776 19880 71780
rect 50296 71836 50360 71840
rect 50296 71780 50300 71836
rect 50300 71780 50356 71836
rect 50356 71780 50360 71836
rect 50296 71776 50360 71780
rect 50376 71836 50440 71840
rect 50376 71780 50380 71836
rect 50380 71780 50436 71836
rect 50436 71780 50440 71836
rect 50376 71776 50440 71780
rect 50456 71836 50520 71840
rect 50456 71780 50460 71836
rect 50460 71780 50516 71836
rect 50516 71780 50520 71836
rect 50456 71776 50520 71780
rect 50536 71836 50600 71840
rect 50536 71780 50540 71836
rect 50540 71780 50596 71836
rect 50596 71780 50600 71836
rect 50536 71776 50600 71780
rect 4216 71292 4280 71296
rect 4216 71236 4220 71292
rect 4220 71236 4276 71292
rect 4276 71236 4280 71292
rect 4216 71232 4280 71236
rect 4296 71292 4360 71296
rect 4296 71236 4300 71292
rect 4300 71236 4356 71292
rect 4356 71236 4360 71292
rect 4296 71232 4360 71236
rect 4376 71292 4440 71296
rect 4376 71236 4380 71292
rect 4380 71236 4436 71292
rect 4436 71236 4440 71292
rect 4376 71232 4440 71236
rect 4456 71292 4520 71296
rect 4456 71236 4460 71292
rect 4460 71236 4516 71292
rect 4516 71236 4520 71292
rect 4456 71232 4520 71236
rect 34936 71292 35000 71296
rect 34936 71236 34940 71292
rect 34940 71236 34996 71292
rect 34996 71236 35000 71292
rect 34936 71232 35000 71236
rect 35016 71292 35080 71296
rect 35016 71236 35020 71292
rect 35020 71236 35076 71292
rect 35076 71236 35080 71292
rect 35016 71232 35080 71236
rect 35096 71292 35160 71296
rect 35096 71236 35100 71292
rect 35100 71236 35156 71292
rect 35156 71236 35160 71292
rect 35096 71232 35160 71236
rect 35176 71292 35240 71296
rect 35176 71236 35180 71292
rect 35180 71236 35236 71292
rect 35236 71236 35240 71292
rect 35176 71232 35240 71236
rect 65656 71292 65720 71296
rect 65656 71236 65660 71292
rect 65660 71236 65716 71292
rect 65716 71236 65720 71292
rect 65656 71232 65720 71236
rect 65736 71292 65800 71296
rect 65736 71236 65740 71292
rect 65740 71236 65796 71292
rect 65796 71236 65800 71292
rect 65736 71232 65800 71236
rect 65816 71292 65880 71296
rect 65816 71236 65820 71292
rect 65820 71236 65876 71292
rect 65876 71236 65880 71292
rect 65816 71232 65880 71236
rect 65896 71292 65960 71296
rect 65896 71236 65900 71292
rect 65900 71236 65956 71292
rect 65956 71236 65960 71292
rect 65896 71232 65960 71236
rect 19576 70748 19640 70752
rect 19576 70692 19580 70748
rect 19580 70692 19636 70748
rect 19636 70692 19640 70748
rect 19576 70688 19640 70692
rect 19656 70748 19720 70752
rect 19656 70692 19660 70748
rect 19660 70692 19716 70748
rect 19716 70692 19720 70748
rect 19656 70688 19720 70692
rect 19736 70748 19800 70752
rect 19736 70692 19740 70748
rect 19740 70692 19796 70748
rect 19796 70692 19800 70748
rect 19736 70688 19800 70692
rect 19816 70748 19880 70752
rect 19816 70692 19820 70748
rect 19820 70692 19876 70748
rect 19876 70692 19880 70748
rect 19816 70688 19880 70692
rect 50296 70748 50360 70752
rect 50296 70692 50300 70748
rect 50300 70692 50356 70748
rect 50356 70692 50360 70748
rect 50296 70688 50360 70692
rect 50376 70748 50440 70752
rect 50376 70692 50380 70748
rect 50380 70692 50436 70748
rect 50436 70692 50440 70748
rect 50376 70688 50440 70692
rect 50456 70748 50520 70752
rect 50456 70692 50460 70748
rect 50460 70692 50516 70748
rect 50516 70692 50520 70748
rect 50456 70688 50520 70692
rect 50536 70748 50600 70752
rect 50536 70692 50540 70748
rect 50540 70692 50596 70748
rect 50596 70692 50600 70748
rect 50536 70688 50600 70692
rect 4216 70204 4280 70208
rect 4216 70148 4220 70204
rect 4220 70148 4276 70204
rect 4276 70148 4280 70204
rect 4216 70144 4280 70148
rect 4296 70204 4360 70208
rect 4296 70148 4300 70204
rect 4300 70148 4356 70204
rect 4356 70148 4360 70204
rect 4296 70144 4360 70148
rect 4376 70204 4440 70208
rect 4376 70148 4380 70204
rect 4380 70148 4436 70204
rect 4436 70148 4440 70204
rect 4376 70144 4440 70148
rect 4456 70204 4520 70208
rect 4456 70148 4460 70204
rect 4460 70148 4516 70204
rect 4516 70148 4520 70204
rect 4456 70144 4520 70148
rect 34936 70204 35000 70208
rect 34936 70148 34940 70204
rect 34940 70148 34996 70204
rect 34996 70148 35000 70204
rect 34936 70144 35000 70148
rect 35016 70204 35080 70208
rect 35016 70148 35020 70204
rect 35020 70148 35076 70204
rect 35076 70148 35080 70204
rect 35016 70144 35080 70148
rect 35096 70204 35160 70208
rect 35096 70148 35100 70204
rect 35100 70148 35156 70204
rect 35156 70148 35160 70204
rect 35096 70144 35160 70148
rect 35176 70204 35240 70208
rect 35176 70148 35180 70204
rect 35180 70148 35236 70204
rect 35236 70148 35240 70204
rect 35176 70144 35240 70148
rect 65656 70204 65720 70208
rect 65656 70148 65660 70204
rect 65660 70148 65716 70204
rect 65716 70148 65720 70204
rect 65656 70144 65720 70148
rect 65736 70204 65800 70208
rect 65736 70148 65740 70204
rect 65740 70148 65796 70204
rect 65796 70148 65800 70204
rect 65736 70144 65800 70148
rect 65816 70204 65880 70208
rect 65816 70148 65820 70204
rect 65820 70148 65876 70204
rect 65876 70148 65880 70204
rect 65816 70144 65880 70148
rect 65896 70204 65960 70208
rect 65896 70148 65900 70204
rect 65900 70148 65956 70204
rect 65956 70148 65960 70204
rect 65896 70144 65960 70148
rect 19576 69660 19640 69664
rect 19576 69604 19580 69660
rect 19580 69604 19636 69660
rect 19636 69604 19640 69660
rect 19576 69600 19640 69604
rect 19656 69660 19720 69664
rect 19656 69604 19660 69660
rect 19660 69604 19716 69660
rect 19716 69604 19720 69660
rect 19656 69600 19720 69604
rect 19736 69660 19800 69664
rect 19736 69604 19740 69660
rect 19740 69604 19796 69660
rect 19796 69604 19800 69660
rect 19736 69600 19800 69604
rect 19816 69660 19880 69664
rect 19816 69604 19820 69660
rect 19820 69604 19876 69660
rect 19876 69604 19880 69660
rect 19816 69600 19880 69604
rect 50296 69660 50360 69664
rect 50296 69604 50300 69660
rect 50300 69604 50356 69660
rect 50356 69604 50360 69660
rect 50296 69600 50360 69604
rect 50376 69660 50440 69664
rect 50376 69604 50380 69660
rect 50380 69604 50436 69660
rect 50436 69604 50440 69660
rect 50376 69600 50440 69604
rect 50456 69660 50520 69664
rect 50456 69604 50460 69660
rect 50460 69604 50516 69660
rect 50516 69604 50520 69660
rect 50456 69600 50520 69604
rect 50536 69660 50600 69664
rect 50536 69604 50540 69660
rect 50540 69604 50596 69660
rect 50596 69604 50600 69660
rect 50536 69600 50600 69604
rect 4216 69116 4280 69120
rect 4216 69060 4220 69116
rect 4220 69060 4276 69116
rect 4276 69060 4280 69116
rect 4216 69056 4280 69060
rect 4296 69116 4360 69120
rect 4296 69060 4300 69116
rect 4300 69060 4356 69116
rect 4356 69060 4360 69116
rect 4296 69056 4360 69060
rect 4376 69116 4440 69120
rect 4376 69060 4380 69116
rect 4380 69060 4436 69116
rect 4436 69060 4440 69116
rect 4376 69056 4440 69060
rect 4456 69116 4520 69120
rect 4456 69060 4460 69116
rect 4460 69060 4516 69116
rect 4516 69060 4520 69116
rect 4456 69056 4520 69060
rect 34936 69116 35000 69120
rect 34936 69060 34940 69116
rect 34940 69060 34996 69116
rect 34996 69060 35000 69116
rect 34936 69056 35000 69060
rect 35016 69116 35080 69120
rect 35016 69060 35020 69116
rect 35020 69060 35076 69116
rect 35076 69060 35080 69116
rect 35016 69056 35080 69060
rect 35096 69116 35160 69120
rect 35096 69060 35100 69116
rect 35100 69060 35156 69116
rect 35156 69060 35160 69116
rect 35096 69056 35160 69060
rect 35176 69116 35240 69120
rect 35176 69060 35180 69116
rect 35180 69060 35236 69116
rect 35236 69060 35240 69116
rect 35176 69056 35240 69060
rect 65656 69116 65720 69120
rect 65656 69060 65660 69116
rect 65660 69060 65716 69116
rect 65716 69060 65720 69116
rect 65656 69056 65720 69060
rect 65736 69116 65800 69120
rect 65736 69060 65740 69116
rect 65740 69060 65796 69116
rect 65796 69060 65800 69116
rect 65736 69056 65800 69060
rect 65816 69116 65880 69120
rect 65816 69060 65820 69116
rect 65820 69060 65876 69116
rect 65876 69060 65880 69116
rect 65816 69056 65880 69060
rect 65896 69116 65960 69120
rect 65896 69060 65900 69116
rect 65900 69060 65956 69116
rect 65956 69060 65960 69116
rect 65896 69056 65960 69060
rect 19576 68572 19640 68576
rect 19576 68516 19580 68572
rect 19580 68516 19636 68572
rect 19636 68516 19640 68572
rect 19576 68512 19640 68516
rect 19656 68572 19720 68576
rect 19656 68516 19660 68572
rect 19660 68516 19716 68572
rect 19716 68516 19720 68572
rect 19656 68512 19720 68516
rect 19736 68572 19800 68576
rect 19736 68516 19740 68572
rect 19740 68516 19796 68572
rect 19796 68516 19800 68572
rect 19736 68512 19800 68516
rect 19816 68572 19880 68576
rect 19816 68516 19820 68572
rect 19820 68516 19876 68572
rect 19876 68516 19880 68572
rect 19816 68512 19880 68516
rect 50296 68572 50360 68576
rect 50296 68516 50300 68572
rect 50300 68516 50356 68572
rect 50356 68516 50360 68572
rect 50296 68512 50360 68516
rect 50376 68572 50440 68576
rect 50376 68516 50380 68572
rect 50380 68516 50436 68572
rect 50436 68516 50440 68572
rect 50376 68512 50440 68516
rect 50456 68572 50520 68576
rect 50456 68516 50460 68572
rect 50460 68516 50516 68572
rect 50516 68516 50520 68572
rect 50456 68512 50520 68516
rect 50536 68572 50600 68576
rect 50536 68516 50540 68572
rect 50540 68516 50596 68572
rect 50596 68516 50600 68572
rect 50536 68512 50600 68516
rect 4216 68028 4280 68032
rect 4216 67972 4220 68028
rect 4220 67972 4276 68028
rect 4276 67972 4280 68028
rect 4216 67968 4280 67972
rect 4296 68028 4360 68032
rect 4296 67972 4300 68028
rect 4300 67972 4356 68028
rect 4356 67972 4360 68028
rect 4296 67968 4360 67972
rect 4376 68028 4440 68032
rect 4376 67972 4380 68028
rect 4380 67972 4436 68028
rect 4436 67972 4440 68028
rect 4376 67968 4440 67972
rect 4456 68028 4520 68032
rect 4456 67972 4460 68028
rect 4460 67972 4516 68028
rect 4516 67972 4520 68028
rect 4456 67968 4520 67972
rect 34936 68028 35000 68032
rect 34936 67972 34940 68028
rect 34940 67972 34996 68028
rect 34996 67972 35000 68028
rect 34936 67968 35000 67972
rect 35016 68028 35080 68032
rect 35016 67972 35020 68028
rect 35020 67972 35076 68028
rect 35076 67972 35080 68028
rect 35016 67968 35080 67972
rect 35096 68028 35160 68032
rect 35096 67972 35100 68028
rect 35100 67972 35156 68028
rect 35156 67972 35160 68028
rect 35096 67968 35160 67972
rect 35176 68028 35240 68032
rect 35176 67972 35180 68028
rect 35180 67972 35236 68028
rect 35236 67972 35240 68028
rect 35176 67968 35240 67972
rect 65656 68028 65720 68032
rect 65656 67972 65660 68028
rect 65660 67972 65716 68028
rect 65716 67972 65720 68028
rect 65656 67968 65720 67972
rect 65736 68028 65800 68032
rect 65736 67972 65740 68028
rect 65740 67972 65796 68028
rect 65796 67972 65800 68028
rect 65736 67968 65800 67972
rect 65816 68028 65880 68032
rect 65816 67972 65820 68028
rect 65820 67972 65876 68028
rect 65876 67972 65880 68028
rect 65816 67968 65880 67972
rect 65896 68028 65960 68032
rect 65896 67972 65900 68028
rect 65900 67972 65956 68028
rect 65956 67972 65960 68028
rect 65896 67968 65960 67972
rect 19576 67484 19640 67488
rect 19576 67428 19580 67484
rect 19580 67428 19636 67484
rect 19636 67428 19640 67484
rect 19576 67424 19640 67428
rect 19656 67484 19720 67488
rect 19656 67428 19660 67484
rect 19660 67428 19716 67484
rect 19716 67428 19720 67484
rect 19656 67424 19720 67428
rect 19736 67484 19800 67488
rect 19736 67428 19740 67484
rect 19740 67428 19796 67484
rect 19796 67428 19800 67484
rect 19736 67424 19800 67428
rect 19816 67484 19880 67488
rect 19816 67428 19820 67484
rect 19820 67428 19876 67484
rect 19876 67428 19880 67484
rect 19816 67424 19880 67428
rect 50296 67484 50360 67488
rect 50296 67428 50300 67484
rect 50300 67428 50356 67484
rect 50356 67428 50360 67484
rect 50296 67424 50360 67428
rect 50376 67484 50440 67488
rect 50376 67428 50380 67484
rect 50380 67428 50436 67484
rect 50436 67428 50440 67484
rect 50376 67424 50440 67428
rect 50456 67484 50520 67488
rect 50456 67428 50460 67484
rect 50460 67428 50516 67484
rect 50516 67428 50520 67484
rect 50456 67424 50520 67428
rect 50536 67484 50600 67488
rect 50536 67428 50540 67484
rect 50540 67428 50596 67484
rect 50596 67428 50600 67484
rect 50536 67424 50600 67428
rect 4216 66940 4280 66944
rect 4216 66884 4220 66940
rect 4220 66884 4276 66940
rect 4276 66884 4280 66940
rect 4216 66880 4280 66884
rect 4296 66940 4360 66944
rect 4296 66884 4300 66940
rect 4300 66884 4356 66940
rect 4356 66884 4360 66940
rect 4296 66880 4360 66884
rect 4376 66940 4440 66944
rect 4376 66884 4380 66940
rect 4380 66884 4436 66940
rect 4436 66884 4440 66940
rect 4376 66880 4440 66884
rect 4456 66940 4520 66944
rect 4456 66884 4460 66940
rect 4460 66884 4516 66940
rect 4516 66884 4520 66940
rect 4456 66880 4520 66884
rect 34936 66940 35000 66944
rect 34936 66884 34940 66940
rect 34940 66884 34996 66940
rect 34996 66884 35000 66940
rect 34936 66880 35000 66884
rect 35016 66940 35080 66944
rect 35016 66884 35020 66940
rect 35020 66884 35076 66940
rect 35076 66884 35080 66940
rect 35016 66880 35080 66884
rect 35096 66940 35160 66944
rect 35096 66884 35100 66940
rect 35100 66884 35156 66940
rect 35156 66884 35160 66940
rect 35096 66880 35160 66884
rect 35176 66940 35240 66944
rect 35176 66884 35180 66940
rect 35180 66884 35236 66940
rect 35236 66884 35240 66940
rect 35176 66880 35240 66884
rect 65656 66940 65720 66944
rect 65656 66884 65660 66940
rect 65660 66884 65716 66940
rect 65716 66884 65720 66940
rect 65656 66880 65720 66884
rect 65736 66940 65800 66944
rect 65736 66884 65740 66940
rect 65740 66884 65796 66940
rect 65796 66884 65800 66940
rect 65736 66880 65800 66884
rect 65816 66940 65880 66944
rect 65816 66884 65820 66940
rect 65820 66884 65876 66940
rect 65876 66884 65880 66940
rect 65816 66880 65880 66884
rect 65896 66940 65960 66944
rect 65896 66884 65900 66940
rect 65900 66884 65956 66940
rect 65956 66884 65960 66940
rect 65896 66880 65960 66884
rect 19576 66396 19640 66400
rect 19576 66340 19580 66396
rect 19580 66340 19636 66396
rect 19636 66340 19640 66396
rect 19576 66336 19640 66340
rect 19656 66396 19720 66400
rect 19656 66340 19660 66396
rect 19660 66340 19716 66396
rect 19716 66340 19720 66396
rect 19656 66336 19720 66340
rect 19736 66396 19800 66400
rect 19736 66340 19740 66396
rect 19740 66340 19796 66396
rect 19796 66340 19800 66396
rect 19736 66336 19800 66340
rect 19816 66396 19880 66400
rect 19816 66340 19820 66396
rect 19820 66340 19876 66396
rect 19876 66340 19880 66396
rect 19816 66336 19880 66340
rect 50296 66396 50360 66400
rect 50296 66340 50300 66396
rect 50300 66340 50356 66396
rect 50356 66340 50360 66396
rect 50296 66336 50360 66340
rect 50376 66396 50440 66400
rect 50376 66340 50380 66396
rect 50380 66340 50436 66396
rect 50436 66340 50440 66396
rect 50376 66336 50440 66340
rect 50456 66396 50520 66400
rect 50456 66340 50460 66396
rect 50460 66340 50516 66396
rect 50516 66340 50520 66396
rect 50456 66336 50520 66340
rect 50536 66396 50600 66400
rect 50536 66340 50540 66396
rect 50540 66340 50596 66396
rect 50596 66340 50600 66396
rect 50536 66336 50600 66340
rect 4216 65852 4280 65856
rect 4216 65796 4220 65852
rect 4220 65796 4276 65852
rect 4276 65796 4280 65852
rect 4216 65792 4280 65796
rect 4296 65852 4360 65856
rect 4296 65796 4300 65852
rect 4300 65796 4356 65852
rect 4356 65796 4360 65852
rect 4296 65792 4360 65796
rect 4376 65852 4440 65856
rect 4376 65796 4380 65852
rect 4380 65796 4436 65852
rect 4436 65796 4440 65852
rect 4376 65792 4440 65796
rect 4456 65852 4520 65856
rect 4456 65796 4460 65852
rect 4460 65796 4516 65852
rect 4516 65796 4520 65852
rect 4456 65792 4520 65796
rect 34936 65852 35000 65856
rect 34936 65796 34940 65852
rect 34940 65796 34996 65852
rect 34996 65796 35000 65852
rect 34936 65792 35000 65796
rect 35016 65852 35080 65856
rect 35016 65796 35020 65852
rect 35020 65796 35076 65852
rect 35076 65796 35080 65852
rect 35016 65792 35080 65796
rect 35096 65852 35160 65856
rect 35096 65796 35100 65852
rect 35100 65796 35156 65852
rect 35156 65796 35160 65852
rect 35096 65792 35160 65796
rect 35176 65852 35240 65856
rect 35176 65796 35180 65852
rect 35180 65796 35236 65852
rect 35236 65796 35240 65852
rect 35176 65792 35240 65796
rect 65656 65852 65720 65856
rect 65656 65796 65660 65852
rect 65660 65796 65716 65852
rect 65716 65796 65720 65852
rect 65656 65792 65720 65796
rect 65736 65852 65800 65856
rect 65736 65796 65740 65852
rect 65740 65796 65796 65852
rect 65796 65796 65800 65852
rect 65736 65792 65800 65796
rect 65816 65852 65880 65856
rect 65816 65796 65820 65852
rect 65820 65796 65876 65852
rect 65876 65796 65880 65852
rect 65816 65792 65880 65796
rect 65896 65852 65960 65856
rect 65896 65796 65900 65852
rect 65900 65796 65956 65852
rect 65956 65796 65960 65852
rect 65896 65792 65960 65796
rect 19576 65308 19640 65312
rect 19576 65252 19580 65308
rect 19580 65252 19636 65308
rect 19636 65252 19640 65308
rect 19576 65248 19640 65252
rect 19656 65308 19720 65312
rect 19656 65252 19660 65308
rect 19660 65252 19716 65308
rect 19716 65252 19720 65308
rect 19656 65248 19720 65252
rect 19736 65308 19800 65312
rect 19736 65252 19740 65308
rect 19740 65252 19796 65308
rect 19796 65252 19800 65308
rect 19736 65248 19800 65252
rect 19816 65308 19880 65312
rect 19816 65252 19820 65308
rect 19820 65252 19876 65308
rect 19876 65252 19880 65308
rect 19816 65248 19880 65252
rect 50296 65308 50360 65312
rect 50296 65252 50300 65308
rect 50300 65252 50356 65308
rect 50356 65252 50360 65308
rect 50296 65248 50360 65252
rect 50376 65308 50440 65312
rect 50376 65252 50380 65308
rect 50380 65252 50436 65308
rect 50436 65252 50440 65308
rect 50376 65248 50440 65252
rect 50456 65308 50520 65312
rect 50456 65252 50460 65308
rect 50460 65252 50516 65308
rect 50516 65252 50520 65308
rect 50456 65248 50520 65252
rect 50536 65308 50600 65312
rect 50536 65252 50540 65308
rect 50540 65252 50596 65308
rect 50596 65252 50600 65308
rect 50536 65248 50600 65252
rect 4216 64764 4280 64768
rect 4216 64708 4220 64764
rect 4220 64708 4276 64764
rect 4276 64708 4280 64764
rect 4216 64704 4280 64708
rect 4296 64764 4360 64768
rect 4296 64708 4300 64764
rect 4300 64708 4356 64764
rect 4356 64708 4360 64764
rect 4296 64704 4360 64708
rect 4376 64764 4440 64768
rect 4376 64708 4380 64764
rect 4380 64708 4436 64764
rect 4436 64708 4440 64764
rect 4376 64704 4440 64708
rect 4456 64764 4520 64768
rect 4456 64708 4460 64764
rect 4460 64708 4516 64764
rect 4516 64708 4520 64764
rect 4456 64704 4520 64708
rect 34936 64764 35000 64768
rect 34936 64708 34940 64764
rect 34940 64708 34996 64764
rect 34996 64708 35000 64764
rect 34936 64704 35000 64708
rect 35016 64764 35080 64768
rect 35016 64708 35020 64764
rect 35020 64708 35076 64764
rect 35076 64708 35080 64764
rect 35016 64704 35080 64708
rect 35096 64764 35160 64768
rect 35096 64708 35100 64764
rect 35100 64708 35156 64764
rect 35156 64708 35160 64764
rect 35096 64704 35160 64708
rect 35176 64764 35240 64768
rect 35176 64708 35180 64764
rect 35180 64708 35236 64764
rect 35236 64708 35240 64764
rect 35176 64704 35240 64708
rect 65656 64764 65720 64768
rect 65656 64708 65660 64764
rect 65660 64708 65716 64764
rect 65716 64708 65720 64764
rect 65656 64704 65720 64708
rect 65736 64764 65800 64768
rect 65736 64708 65740 64764
rect 65740 64708 65796 64764
rect 65796 64708 65800 64764
rect 65736 64704 65800 64708
rect 65816 64764 65880 64768
rect 65816 64708 65820 64764
rect 65820 64708 65876 64764
rect 65876 64708 65880 64764
rect 65816 64704 65880 64708
rect 65896 64764 65960 64768
rect 65896 64708 65900 64764
rect 65900 64708 65956 64764
rect 65956 64708 65960 64764
rect 65896 64704 65960 64708
rect 19576 64220 19640 64224
rect 19576 64164 19580 64220
rect 19580 64164 19636 64220
rect 19636 64164 19640 64220
rect 19576 64160 19640 64164
rect 19656 64220 19720 64224
rect 19656 64164 19660 64220
rect 19660 64164 19716 64220
rect 19716 64164 19720 64220
rect 19656 64160 19720 64164
rect 19736 64220 19800 64224
rect 19736 64164 19740 64220
rect 19740 64164 19796 64220
rect 19796 64164 19800 64220
rect 19736 64160 19800 64164
rect 19816 64220 19880 64224
rect 19816 64164 19820 64220
rect 19820 64164 19876 64220
rect 19876 64164 19880 64220
rect 19816 64160 19880 64164
rect 50296 64220 50360 64224
rect 50296 64164 50300 64220
rect 50300 64164 50356 64220
rect 50356 64164 50360 64220
rect 50296 64160 50360 64164
rect 50376 64220 50440 64224
rect 50376 64164 50380 64220
rect 50380 64164 50436 64220
rect 50436 64164 50440 64220
rect 50376 64160 50440 64164
rect 50456 64220 50520 64224
rect 50456 64164 50460 64220
rect 50460 64164 50516 64220
rect 50516 64164 50520 64220
rect 50456 64160 50520 64164
rect 50536 64220 50600 64224
rect 50536 64164 50540 64220
rect 50540 64164 50596 64220
rect 50596 64164 50600 64220
rect 50536 64160 50600 64164
rect 4216 63676 4280 63680
rect 4216 63620 4220 63676
rect 4220 63620 4276 63676
rect 4276 63620 4280 63676
rect 4216 63616 4280 63620
rect 4296 63676 4360 63680
rect 4296 63620 4300 63676
rect 4300 63620 4356 63676
rect 4356 63620 4360 63676
rect 4296 63616 4360 63620
rect 4376 63676 4440 63680
rect 4376 63620 4380 63676
rect 4380 63620 4436 63676
rect 4436 63620 4440 63676
rect 4376 63616 4440 63620
rect 4456 63676 4520 63680
rect 4456 63620 4460 63676
rect 4460 63620 4516 63676
rect 4516 63620 4520 63676
rect 4456 63616 4520 63620
rect 34936 63676 35000 63680
rect 34936 63620 34940 63676
rect 34940 63620 34996 63676
rect 34996 63620 35000 63676
rect 34936 63616 35000 63620
rect 35016 63676 35080 63680
rect 35016 63620 35020 63676
rect 35020 63620 35076 63676
rect 35076 63620 35080 63676
rect 35016 63616 35080 63620
rect 35096 63676 35160 63680
rect 35096 63620 35100 63676
rect 35100 63620 35156 63676
rect 35156 63620 35160 63676
rect 35096 63616 35160 63620
rect 35176 63676 35240 63680
rect 35176 63620 35180 63676
rect 35180 63620 35236 63676
rect 35236 63620 35240 63676
rect 35176 63616 35240 63620
rect 65656 63676 65720 63680
rect 65656 63620 65660 63676
rect 65660 63620 65716 63676
rect 65716 63620 65720 63676
rect 65656 63616 65720 63620
rect 65736 63676 65800 63680
rect 65736 63620 65740 63676
rect 65740 63620 65796 63676
rect 65796 63620 65800 63676
rect 65736 63616 65800 63620
rect 65816 63676 65880 63680
rect 65816 63620 65820 63676
rect 65820 63620 65876 63676
rect 65876 63620 65880 63676
rect 65816 63616 65880 63620
rect 65896 63676 65960 63680
rect 65896 63620 65900 63676
rect 65900 63620 65956 63676
rect 65956 63620 65960 63676
rect 65896 63616 65960 63620
rect 19576 63132 19640 63136
rect 19576 63076 19580 63132
rect 19580 63076 19636 63132
rect 19636 63076 19640 63132
rect 19576 63072 19640 63076
rect 19656 63132 19720 63136
rect 19656 63076 19660 63132
rect 19660 63076 19716 63132
rect 19716 63076 19720 63132
rect 19656 63072 19720 63076
rect 19736 63132 19800 63136
rect 19736 63076 19740 63132
rect 19740 63076 19796 63132
rect 19796 63076 19800 63132
rect 19736 63072 19800 63076
rect 19816 63132 19880 63136
rect 19816 63076 19820 63132
rect 19820 63076 19876 63132
rect 19876 63076 19880 63132
rect 19816 63072 19880 63076
rect 50296 63132 50360 63136
rect 50296 63076 50300 63132
rect 50300 63076 50356 63132
rect 50356 63076 50360 63132
rect 50296 63072 50360 63076
rect 50376 63132 50440 63136
rect 50376 63076 50380 63132
rect 50380 63076 50436 63132
rect 50436 63076 50440 63132
rect 50376 63072 50440 63076
rect 50456 63132 50520 63136
rect 50456 63076 50460 63132
rect 50460 63076 50516 63132
rect 50516 63076 50520 63132
rect 50456 63072 50520 63076
rect 50536 63132 50600 63136
rect 50536 63076 50540 63132
rect 50540 63076 50596 63132
rect 50596 63076 50600 63132
rect 50536 63072 50600 63076
rect 4216 62588 4280 62592
rect 4216 62532 4220 62588
rect 4220 62532 4276 62588
rect 4276 62532 4280 62588
rect 4216 62528 4280 62532
rect 4296 62588 4360 62592
rect 4296 62532 4300 62588
rect 4300 62532 4356 62588
rect 4356 62532 4360 62588
rect 4296 62528 4360 62532
rect 4376 62588 4440 62592
rect 4376 62532 4380 62588
rect 4380 62532 4436 62588
rect 4436 62532 4440 62588
rect 4376 62528 4440 62532
rect 4456 62588 4520 62592
rect 4456 62532 4460 62588
rect 4460 62532 4516 62588
rect 4516 62532 4520 62588
rect 4456 62528 4520 62532
rect 34936 62588 35000 62592
rect 34936 62532 34940 62588
rect 34940 62532 34996 62588
rect 34996 62532 35000 62588
rect 34936 62528 35000 62532
rect 35016 62588 35080 62592
rect 35016 62532 35020 62588
rect 35020 62532 35076 62588
rect 35076 62532 35080 62588
rect 35016 62528 35080 62532
rect 35096 62588 35160 62592
rect 35096 62532 35100 62588
rect 35100 62532 35156 62588
rect 35156 62532 35160 62588
rect 35096 62528 35160 62532
rect 35176 62588 35240 62592
rect 35176 62532 35180 62588
rect 35180 62532 35236 62588
rect 35236 62532 35240 62588
rect 35176 62528 35240 62532
rect 65656 62588 65720 62592
rect 65656 62532 65660 62588
rect 65660 62532 65716 62588
rect 65716 62532 65720 62588
rect 65656 62528 65720 62532
rect 65736 62588 65800 62592
rect 65736 62532 65740 62588
rect 65740 62532 65796 62588
rect 65796 62532 65800 62588
rect 65736 62528 65800 62532
rect 65816 62588 65880 62592
rect 65816 62532 65820 62588
rect 65820 62532 65876 62588
rect 65876 62532 65880 62588
rect 65816 62528 65880 62532
rect 65896 62588 65960 62592
rect 65896 62532 65900 62588
rect 65900 62532 65956 62588
rect 65956 62532 65960 62588
rect 65896 62528 65960 62532
rect 19576 62044 19640 62048
rect 19576 61988 19580 62044
rect 19580 61988 19636 62044
rect 19636 61988 19640 62044
rect 19576 61984 19640 61988
rect 19656 62044 19720 62048
rect 19656 61988 19660 62044
rect 19660 61988 19716 62044
rect 19716 61988 19720 62044
rect 19656 61984 19720 61988
rect 19736 62044 19800 62048
rect 19736 61988 19740 62044
rect 19740 61988 19796 62044
rect 19796 61988 19800 62044
rect 19736 61984 19800 61988
rect 19816 62044 19880 62048
rect 19816 61988 19820 62044
rect 19820 61988 19876 62044
rect 19876 61988 19880 62044
rect 19816 61984 19880 61988
rect 50296 62044 50360 62048
rect 50296 61988 50300 62044
rect 50300 61988 50356 62044
rect 50356 61988 50360 62044
rect 50296 61984 50360 61988
rect 50376 62044 50440 62048
rect 50376 61988 50380 62044
rect 50380 61988 50436 62044
rect 50436 61988 50440 62044
rect 50376 61984 50440 61988
rect 50456 62044 50520 62048
rect 50456 61988 50460 62044
rect 50460 61988 50516 62044
rect 50516 61988 50520 62044
rect 50456 61984 50520 61988
rect 50536 62044 50600 62048
rect 50536 61988 50540 62044
rect 50540 61988 50596 62044
rect 50596 61988 50600 62044
rect 50536 61984 50600 61988
rect 4216 61500 4280 61504
rect 4216 61444 4220 61500
rect 4220 61444 4276 61500
rect 4276 61444 4280 61500
rect 4216 61440 4280 61444
rect 4296 61500 4360 61504
rect 4296 61444 4300 61500
rect 4300 61444 4356 61500
rect 4356 61444 4360 61500
rect 4296 61440 4360 61444
rect 4376 61500 4440 61504
rect 4376 61444 4380 61500
rect 4380 61444 4436 61500
rect 4436 61444 4440 61500
rect 4376 61440 4440 61444
rect 4456 61500 4520 61504
rect 4456 61444 4460 61500
rect 4460 61444 4516 61500
rect 4516 61444 4520 61500
rect 4456 61440 4520 61444
rect 34936 61500 35000 61504
rect 34936 61444 34940 61500
rect 34940 61444 34996 61500
rect 34996 61444 35000 61500
rect 34936 61440 35000 61444
rect 35016 61500 35080 61504
rect 35016 61444 35020 61500
rect 35020 61444 35076 61500
rect 35076 61444 35080 61500
rect 35016 61440 35080 61444
rect 35096 61500 35160 61504
rect 35096 61444 35100 61500
rect 35100 61444 35156 61500
rect 35156 61444 35160 61500
rect 35096 61440 35160 61444
rect 35176 61500 35240 61504
rect 35176 61444 35180 61500
rect 35180 61444 35236 61500
rect 35236 61444 35240 61500
rect 35176 61440 35240 61444
rect 65656 61500 65720 61504
rect 65656 61444 65660 61500
rect 65660 61444 65716 61500
rect 65716 61444 65720 61500
rect 65656 61440 65720 61444
rect 65736 61500 65800 61504
rect 65736 61444 65740 61500
rect 65740 61444 65796 61500
rect 65796 61444 65800 61500
rect 65736 61440 65800 61444
rect 65816 61500 65880 61504
rect 65816 61444 65820 61500
rect 65820 61444 65876 61500
rect 65876 61444 65880 61500
rect 65816 61440 65880 61444
rect 65896 61500 65960 61504
rect 65896 61444 65900 61500
rect 65900 61444 65956 61500
rect 65956 61444 65960 61500
rect 65896 61440 65960 61444
rect 19576 60956 19640 60960
rect 19576 60900 19580 60956
rect 19580 60900 19636 60956
rect 19636 60900 19640 60956
rect 19576 60896 19640 60900
rect 19656 60956 19720 60960
rect 19656 60900 19660 60956
rect 19660 60900 19716 60956
rect 19716 60900 19720 60956
rect 19656 60896 19720 60900
rect 19736 60956 19800 60960
rect 19736 60900 19740 60956
rect 19740 60900 19796 60956
rect 19796 60900 19800 60956
rect 19736 60896 19800 60900
rect 19816 60956 19880 60960
rect 19816 60900 19820 60956
rect 19820 60900 19876 60956
rect 19876 60900 19880 60956
rect 19816 60896 19880 60900
rect 50296 60956 50360 60960
rect 50296 60900 50300 60956
rect 50300 60900 50356 60956
rect 50356 60900 50360 60956
rect 50296 60896 50360 60900
rect 50376 60956 50440 60960
rect 50376 60900 50380 60956
rect 50380 60900 50436 60956
rect 50436 60900 50440 60956
rect 50376 60896 50440 60900
rect 50456 60956 50520 60960
rect 50456 60900 50460 60956
rect 50460 60900 50516 60956
rect 50516 60900 50520 60956
rect 50456 60896 50520 60900
rect 50536 60956 50600 60960
rect 50536 60900 50540 60956
rect 50540 60900 50596 60956
rect 50596 60900 50600 60956
rect 50536 60896 50600 60900
rect 4216 60412 4280 60416
rect 4216 60356 4220 60412
rect 4220 60356 4276 60412
rect 4276 60356 4280 60412
rect 4216 60352 4280 60356
rect 4296 60412 4360 60416
rect 4296 60356 4300 60412
rect 4300 60356 4356 60412
rect 4356 60356 4360 60412
rect 4296 60352 4360 60356
rect 4376 60412 4440 60416
rect 4376 60356 4380 60412
rect 4380 60356 4436 60412
rect 4436 60356 4440 60412
rect 4376 60352 4440 60356
rect 4456 60412 4520 60416
rect 4456 60356 4460 60412
rect 4460 60356 4516 60412
rect 4516 60356 4520 60412
rect 4456 60352 4520 60356
rect 34936 60412 35000 60416
rect 34936 60356 34940 60412
rect 34940 60356 34996 60412
rect 34996 60356 35000 60412
rect 34936 60352 35000 60356
rect 35016 60412 35080 60416
rect 35016 60356 35020 60412
rect 35020 60356 35076 60412
rect 35076 60356 35080 60412
rect 35016 60352 35080 60356
rect 35096 60412 35160 60416
rect 35096 60356 35100 60412
rect 35100 60356 35156 60412
rect 35156 60356 35160 60412
rect 35096 60352 35160 60356
rect 35176 60412 35240 60416
rect 35176 60356 35180 60412
rect 35180 60356 35236 60412
rect 35236 60356 35240 60412
rect 35176 60352 35240 60356
rect 65656 60412 65720 60416
rect 65656 60356 65660 60412
rect 65660 60356 65716 60412
rect 65716 60356 65720 60412
rect 65656 60352 65720 60356
rect 65736 60412 65800 60416
rect 65736 60356 65740 60412
rect 65740 60356 65796 60412
rect 65796 60356 65800 60412
rect 65736 60352 65800 60356
rect 65816 60412 65880 60416
rect 65816 60356 65820 60412
rect 65820 60356 65876 60412
rect 65876 60356 65880 60412
rect 65816 60352 65880 60356
rect 65896 60412 65960 60416
rect 65896 60356 65900 60412
rect 65900 60356 65956 60412
rect 65956 60356 65960 60412
rect 65896 60352 65960 60356
rect 19576 59868 19640 59872
rect 19576 59812 19580 59868
rect 19580 59812 19636 59868
rect 19636 59812 19640 59868
rect 19576 59808 19640 59812
rect 19656 59868 19720 59872
rect 19656 59812 19660 59868
rect 19660 59812 19716 59868
rect 19716 59812 19720 59868
rect 19656 59808 19720 59812
rect 19736 59868 19800 59872
rect 19736 59812 19740 59868
rect 19740 59812 19796 59868
rect 19796 59812 19800 59868
rect 19736 59808 19800 59812
rect 19816 59868 19880 59872
rect 19816 59812 19820 59868
rect 19820 59812 19876 59868
rect 19876 59812 19880 59868
rect 19816 59808 19880 59812
rect 50296 59868 50360 59872
rect 50296 59812 50300 59868
rect 50300 59812 50356 59868
rect 50356 59812 50360 59868
rect 50296 59808 50360 59812
rect 50376 59868 50440 59872
rect 50376 59812 50380 59868
rect 50380 59812 50436 59868
rect 50436 59812 50440 59868
rect 50376 59808 50440 59812
rect 50456 59868 50520 59872
rect 50456 59812 50460 59868
rect 50460 59812 50516 59868
rect 50516 59812 50520 59868
rect 50456 59808 50520 59812
rect 50536 59868 50600 59872
rect 50536 59812 50540 59868
rect 50540 59812 50596 59868
rect 50596 59812 50600 59868
rect 50536 59808 50600 59812
rect 4216 59324 4280 59328
rect 4216 59268 4220 59324
rect 4220 59268 4276 59324
rect 4276 59268 4280 59324
rect 4216 59264 4280 59268
rect 4296 59324 4360 59328
rect 4296 59268 4300 59324
rect 4300 59268 4356 59324
rect 4356 59268 4360 59324
rect 4296 59264 4360 59268
rect 4376 59324 4440 59328
rect 4376 59268 4380 59324
rect 4380 59268 4436 59324
rect 4436 59268 4440 59324
rect 4376 59264 4440 59268
rect 4456 59324 4520 59328
rect 4456 59268 4460 59324
rect 4460 59268 4516 59324
rect 4516 59268 4520 59324
rect 4456 59264 4520 59268
rect 34936 59324 35000 59328
rect 34936 59268 34940 59324
rect 34940 59268 34996 59324
rect 34996 59268 35000 59324
rect 34936 59264 35000 59268
rect 35016 59324 35080 59328
rect 35016 59268 35020 59324
rect 35020 59268 35076 59324
rect 35076 59268 35080 59324
rect 35016 59264 35080 59268
rect 35096 59324 35160 59328
rect 35096 59268 35100 59324
rect 35100 59268 35156 59324
rect 35156 59268 35160 59324
rect 35096 59264 35160 59268
rect 35176 59324 35240 59328
rect 35176 59268 35180 59324
rect 35180 59268 35236 59324
rect 35236 59268 35240 59324
rect 35176 59264 35240 59268
rect 65656 59324 65720 59328
rect 65656 59268 65660 59324
rect 65660 59268 65716 59324
rect 65716 59268 65720 59324
rect 65656 59264 65720 59268
rect 65736 59324 65800 59328
rect 65736 59268 65740 59324
rect 65740 59268 65796 59324
rect 65796 59268 65800 59324
rect 65736 59264 65800 59268
rect 65816 59324 65880 59328
rect 65816 59268 65820 59324
rect 65820 59268 65876 59324
rect 65876 59268 65880 59324
rect 65816 59264 65880 59268
rect 65896 59324 65960 59328
rect 65896 59268 65900 59324
rect 65900 59268 65956 59324
rect 65956 59268 65960 59324
rect 65896 59264 65960 59268
rect 19576 58780 19640 58784
rect 19576 58724 19580 58780
rect 19580 58724 19636 58780
rect 19636 58724 19640 58780
rect 19576 58720 19640 58724
rect 19656 58780 19720 58784
rect 19656 58724 19660 58780
rect 19660 58724 19716 58780
rect 19716 58724 19720 58780
rect 19656 58720 19720 58724
rect 19736 58780 19800 58784
rect 19736 58724 19740 58780
rect 19740 58724 19796 58780
rect 19796 58724 19800 58780
rect 19736 58720 19800 58724
rect 19816 58780 19880 58784
rect 19816 58724 19820 58780
rect 19820 58724 19876 58780
rect 19876 58724 19880 58780
rect 19816 58720 19880 58724
rect 50296 58780 50360 58784
rect 50296 58724 50300 58780
rect 50300 58724 50356 58780
rect 50356 58724 50360 58780
rect 50296 58720 50360 58724
rect 50376 58780 50440 58784
rect 50376 58724 50380 58780
rect 50380 58724 50436 58780
rect 50436 58724 50440 58780
rect 50376 58720 50440 58724
rect 50456 58780 50520 58784
rect 50456 58724 50460 58780
rect 50460 58724 50516 58780
rect 50516 58724 50520 58780
rect 50456 58720 50520 58724
rect 50536 58780 50600 58784
rect 50536 58724 50540 58780
rect 50540 58724 50596 58780
rect 50596 58724 50600 58780
rect 50536 58720 50600 58724
rect 4216 58236 4280 58240
rect 4216 58180 4220 58236
rect 4220 58180 4276 58236
rect 4276 58180 4280 58236
rect 4216 58176 4280 58180
rect 4296 58236 4360 58240
rect 4296 58180 4300 58236
rect 4300 58180 4356 58236
rect 4356 58180 4360 58236
rect 4296 58176 4360 58180
rect 4376 58236 4440 58240
rect 4376 58180 4380 58236
rect 4380 58180 4436 58236
rect 4436 58180 4440 58236
rect 4376 58176 4440 58180
rect 4456 58236 4520 58240
rect 4456 58180 4460 58236
rect 4460 58180 4516 58236
rect 4516 58180 4520 58236
rect 4456 58176 4520 58180
rect 34936 58236 35000 58240
rect 34936 58180 34940 58236
rect 34940 58180 34996 58236
rect 34996 58180 35000 58236
rect 34936 58176 35000 58180
rect 35016 58236 35080 58240
rect 35016 58180 35020 58236
rect 35020 58180 35076 58236
rect 35076 58180 35080 58236
rect 35016 58176 35080 58180
rect 35096 58236 35160 58240
rect 35096 58180 35100 58236
rect 35100 58180 35156 58236
rect 35156 58180 35160 58236
rect 35096 58176 35160 58180
rect 35176 58236 35240 58240
rect 35176 58180 35180 58236
rect 35180 58180 35236 58236
rect 35236 58180 35240 58236
rect 35176 58176 35240 58180
rect 65656 58236 65720 58240
rect 65656 58180 65660 58236
rect 65660 58180 65716 58236
rect 65716 58180 65720 58236
rect 65656 58176 65720 58180
rect 65736 58236 65800 58240
rect 65736 58180 65740 58236
rect 65740 58180 65796 58236
rect 65796 58180 65800 58236
rect 65736 58176 65800 58180
rect 65816 58236 65880 58240
rect 65816 58180 65820 58236
rect 65820 58180 65876 58236
rect 65876 58180 65880 58236
rect 65816 58176 65880 58180
rect 65896 58236 65960 58240
rect 65896 58180 65900 58236
rect 65900 58180 65956 58236
rect 65956 58180 65960 58236
rect 65896 58176 65960 58180
rect 19576 57692 19640 57696
rect 19576 57636 19580 57692
rect 19580 57636 19636 57692
rect 19636 57636 19640 57692
rect 19576 57632 19640 57636
rect 19656 57692 19720 57696
rect 19656 57636 19660 57692
rect 19660 57636 19716 57692
rect 19716 57636 19720 57692
rect 19656 57632 19720 57636
rect 19736 57692 19800 57696
rect 19736 57636 19740 57692
rect 19740 57636 19796 57692
rect 19796 57636 19800 57692
rect 19736 57632 19800 57636
rect 19816 57692 19880 57696
rect 19816 57636 19820 57692
rect 19820 57636 19876 57692
rect 19876 57636 19880 57692
rect 19816 57632 19880 57636
rect 50296 57692 50360 57696
rect 50296 57636 50300 57692
rect 50300 57636 50356 57692
rect 50356 57636 50360 57692
rect 50296 57632 50360 57636
rect 50376 57692 50440 57696
rect 50376 57636 50380 57692
rect 50380 57636 50436 57692
rect 50436 57636 50440 57692
rect 50376 57632 50440 57636
rect 50456 57692 50520 57696
rect 50456 57636 50460 57692
rect 50460 57636 50516 57692
rect 50516 57636 50520 57692
rect 50456 57632 50520 57636
rect 50536 57692 50600 57696
rect 50536 57636 50540 57692
rect 50540 57636 50596 57692
rect 50596 57636 50600 57692
rect 50536 57632 50600 57636
rect 4216 57148 4280 57152
rect 4216 57092 4220 57148
rect 4220 57092 4276 57148
rect 4276 57092 4280 57148
rect 4216 57088 4280 57092
rect 4296 57148 4360 57152
rect 4296 57092 4300 57148
rect 4300 57092 4356 57148
rect 4356 57092 4360 57148
rect 4296 57088 4360 57092
rect 4376 57148 4440 57152
rect 4376 57092 4380 57148
rect 4380 57092 4436 57148
rect 4436 57092 4440 57148
rect 4376 57088 4440 57092
rect 4456 57148 4520 57152
rect 4456 57092 4460 57148
rect 4460 57092 4516 57148
rect 4516 57092 4520 57148
rect 4456 57088 4520 57092
rect 34936 57148 35000 57152
rect 34936 57092 34940 57148
rect 34940 57092 34996 57148
rect 34996 57092 35000 57148
rect 34936 57088 35000 57092
rect 35016 57148 35080 57152
rect 35016 57092 35020 57148
rect 35020 57092 35076 57148
rect 35076 57092 35080 57148
rect 35016 57088 35080 57092
rect 35096 57148 35160 57152
rect 35096 57092 35100 57148
rect 35100 57092 35156 57148
rect 35156 57092 35160 57148
rect 35096 57088 35160 57092
rect 35176 57148 35240 57152
rect 35176 57092 35180 57148
rect 35180 57092 35236 57148
rect 35236 57092 35240 57148
rect 35176 57088 35240 57092
rect 65656 57148 65720 57152
rect 65656 57092 65660 57148
rect 65660 57092 65716 57148
rect 65716 57092 65720 57148
rect 65656 57088 65720 57092
rect 65736 57148 65800 57152
rect 65736 57092 65740 57148
rect 65740 57092 65796 57148
rect 65796 57092 65800 57148
rect 65736 57088 65800 57092
rect 65816 57148 65880 57152
rect 65816 57092 65820 57148
rect 65820 57092 65876 57148
rect 65876 57092 65880 57148
rect 65816 57088 65880 57092
rect 65896 57148 65960 57152
rect 65896 57092 65900 57148
rect 65900 57092 65956 57148
rect 65956 57092 65960 57148
rect 65896 57088 65960 57092
rect 19576 56604 19640 56608
rect 19576 56548 19580 56604
rect 19580 56548 19636 56604
rect 19636 56548 19640 56604
rect 19576 56544 19640 56548
rect 19656 56604 19720 56608
rect 19656 56548 19660 56604
rect 19660 56548 19716 56604
rect 19716 56548 19720 56604
rect 19656 56544 19720 56548
rect 19736 56604 19800 56608
rect 19736 56548 19740 56604
rect 19740 56548 19796 56604
rect 19796 56548 19800 56604
rect 19736 56544 19800 56548
rect 19816 56604 19880 56608
rect 19816 56548 19820 56604
rect 19820 56548 19876 56604
rect 19876 56548 19880 56604
rect 19816 56544 19880 56548
rect 50296 56604 50360 56608
rect 50296 56548 50300 56604
rect 50300 56548 50356 56604
rect 50356 56548 50360 56604
rect 50296 56544 50360 56548
rect 50376 56604 50440 56608
rect 50376 56548 50380 56604
rect 50380 56548 50436 56604
rect 50436 56548 50440 56604
rect 50376 56544 50440 56548
rect 50456 56604 50520 56608
rect 50456 56548 50460 56604
rect 50460 56548 50516 56604
rect 50516 56548 50520 56604
rect 50456 56544 50520 56548
rect 50536 56604 50600 56608
rect 50536 56548 50540 56604
rect 50540 56548 50596 56604
rect 50596 56548 50600 56604
rect 50536 56544 50600 56548
rect 4216 56060 4280 56064
rect 4216 56004 4220 56060
rect 4220 56004 4276 56060
rect 4276 56004 4280 56060
rect 4216 56000 4280 56004
rect 4296 56060 4360 56064
rect 4296 56004 4300 56060
rect 4300 56004 4356 56060
rect 4356 56004 4360 56060
rect 4296 56000 4360 56004
rect 4376 56060 4440 56064
rect 4376 56004 4380 56060
rect 4380 56004 4436 56060
rect 4436 56004 4440 56060
rect 4376 56000 4440 56004
rect 4456 56060 4520 56064
rect 4456 56004 4460 56060
rect 4460 56004 4516 56060
rect 4516 56004 4520 56060
rect 4456 56000 4520 56004
rect 34936 56060 35000 56064
rect 34936 56004 34940 56060
rect 34940 56004 34996 56060
rect 34996 56004 35000 56060
rect 34936 56000 35000 56004
rect 35016 56060 35080 56064
rect 35016 56004 35020 56060
rect 35020 56004 35076 56060
rect 35076 56004 35080 56060
rect 35016 56000 35080 56004
rect 35096 56060 35160 56064
rect 35096 56004 35100 56060
rect 35100 56004 35156 56060
rect 35156 56004 35160 56060
rect 35096 56000 35160 56004
rect 35176 56060 35240 56064
rect 35176 56004 35180 56060
rect 35180 56004 35236 56060
rect 35236 56004 35240 56060
rect 35176 56000 35240 56004
rect 65656 56060 65720 56064
rect 65656 56004 65660 56060
rect 65660 56004 65716 56060
rect 65716 56004 65720 56060
rect 65656 56000 65720 56004
rect 65736 56060 65800 56064
rect 65736 56004 65740 56060
rect 65740 56004 65796 56060
rect 65796 56004 65800 56060
rect 65736 56000 65800 56004
rect 65816 56060 65880 56064
rect 65816 56004 65820 56060
rect 65820 56004 65876 56060
rect 65876 56004 65880 56060
rect 65816 56000 65880 56004
rect 65896 56060 65960 56064
rect 65896 56004 65900 56060
rect 65900 56004 65956 56060
rect 65956 56004 65960 56060
rect 65896 56000 65960 56004
rect 19576 55516 19640 55520
rect 19576 55460 19580 55516
rect 19580 55460 19636 55516
rect 19636 55460 19640 55516
rect 19576 55456 19640 55460
rect 19656 55516 19720 55520
rect 19656 55460 19660 55516
rect 19660 55460 19716 55516
rect 19716 55460 19720 55516
rect 19656 55456 19720 55460
rect 19736 55516 19800 55520
rect 19736 55460 19740 55516
rect 19740 55460 19796 55516
rect 19796 55460 19800 55516
rect 19736 55456 19800 55460
rect 19816 55516 19880 55520
rect 19816 55460 19820 55516
rect 19820 55460 19876 55516
rect 19876 55460 19880 55516
rect 19816 55456 19880 55460
rect 50296 55516 50360 55520
rect 50296 55460 50300 55516
rect 50300 55460 50356 55516
rect 50356 55460 50360 55516
rect 50296 55456 50360 55460
rect 50376 55516 50440 55520
rect 50376 55460 50380 55516
rect 50380 55460 50436 55516
rect 50436 55460 50440 55516
rect 50376 55456 50440 55460
rect 50456 55516 50520 55520
rect 50456 55460 50460 55516
rect 50460 55460 50516 55516
rect 50516 55460 50520 55516
rect 50456 55456 50520 55460
rect 50536 55516 50600 55520
rect 50536 55460 50540 55516
rect 50540 55460 50596 55516
rect 50596 55460 50600 55516
rect 50536 55456 50600 55460
rect 4216 54972 4280 54976
rect 4216 54916 4220 54972
rect 4220 54916 4276 54972
rect 4276 54916 4280 54972
rect 4216 54912 4280 54916
rect 4296 54972 4360 54976
rect 4296 54916 4300 54972
rect 4300 54916 4356 54972
rect 4356 54916 4360 54972
rect 4296 54912 4360 54916
rect 4376 54972 4440 54976
rect 4376 54916 4380 54972
rect 4380 54916 4436 54972
rect 4436 54916 4440 54972
rect 4376 54912 4440 54916
rect 4456 54972 4520 54976
rect 4456 54916 4460 54972
rect 4460 54916 4516 54972
rect 4516 54916 4520 54972
rect 4456 54912 4520 54916
rect 34936 54972 35000 54976
rect 34936 54916 34940 54972
rect 34940 54916 34996 54972
rect 34996 54916 35000 54972
rect 34936 54912 35000 54916
rect 35016 54972 35080 54976
rect 35016 54916 35020 54972
rect 35020 54916 35076 54972
rect 35076 54916 35080 54972
rect 35016 54912 35080 54916
rect 35096 54972 35160 54976
rect 35096 54916 35100 54972
rect 35100 54916 35156 54972
rect 35156 54916 35160 54972
rect 35096 54912 35160 54916
rect 35176 54972 35240 54976
rect 35176 54916 35180 54972
rect 35180 54916 35236 54972
rect 35236 54916 35240 54972
rect 35176 54912 35240 54916
rect 65656 54972 65720 54976
rect 65656 54916 65660 54972
rect 65660 54916 65716 54972
rect 65716 54916 65720 54972
rect 65656 54912 65720 54916
rect 65736 54972 65800 54976
rect 65736 54916 65740 54972
rect 65740 54916 65796 54972
rect 65796 54916 65800 54972
rect 65736 54912 65800 54916
rect 65816 54972 65880 54976
rect 65816 54916 65820 54972
rect 65820 54916 65876 54972
rect 65876 54916 65880 54972
rect 65816 54912 65880 54916
rect 65896 54972 65960 54976
rect 65896 54916 65900 54972
rect 65900 54916 65956 54972
rect 65956 54916 65960 54972
rect 65896 54912 65960 54916
rect 19576 54428 19640 54432
rect 19576 54372 19580 54428
rect 19580 54372 19636 54428
rect 19636 54372 19640 54428
rect 19576 54368 19640 54372
rect 19656 54428 19720 54432
rect 19656 54372 19660 54428
rect 19660 54372 19716 54428
rect 19716 54372 19720 54428
rect 19656 54368 19720 54372
rect 19736 54428 19800 54432
rect 19736 54372 19740 54428
rect 19740 54372 19796 54428
rect 19796 54372 19800 54428
rect 19736 54368 19800 54372
rect 19816 54428 19880 54432
rect 19816 54372 19820 54428
rect 19820 54372 19876 54428
rect 19876 54372 19880 54428
rect 19816 54368 19880 54372
rect 50296 54428 50360 54432
rect 50296 54372 50300 54428
rect 50300 54372 50356 54428
rect 50356 54372 50360 54428
rect 50296 54368 50360 54372
rect 50376 54428 50440 54432
rect 50376 54372 50380 54428
rect 50380 54372 50436 54428
rect 50436 54372 50440 54428
rect 50376 54368 50440 54372
rect 50456 54428 50520 54432
rect 50456 54372 50460 54428
rect 50460 54372 50516 54428
rect 50516 54372 50520 54428
rect 50456 54368 50520 54372
rect 50536 54428 50600 54432
rect 50536 54372 50540 54428
rect 50540 54372 50596 54428
rect 50596 54372 50600 54428
rect 50536 54368 50600 54372
rect 4216 53884 4280 53888
rect 4216 53828 4220 53884
rect 4220 53828 4276 53884
rect 4276 53828 4280 53884
rect 4216 53824 4280 53828
rect 4296 53884 4360 53888
rect 4296 53828 4300 53884
rect 4300 53828 4356 53884
rect 4356 53828 4360 53884
rect 4296 53824 4360 53828
rect 4376 53884 4440 53888
rect 4376 53828 4380 53884
rect 4380 53828 4436 53884
rect 4436 53828 4440 53884
rect 4376 53824 4440 53828
rect 4456 53884 4520 53888
rect 4456 53828 4460 53884
rect 4460 53828 4516 53884
rect 4516 53828 4520 53884
rect 4456 53824 4520 53828
rect 34936 53884 35000 53888
rect 34936 53828 34940 53884
rect 34940 53828 34996 53884
rect 34996 53828 35000 53884
rect 34936 53824 35000 53828
rect 35016 53884 35080 53888
rect 35016 53828 35020 53884
rect 35020 53828 35076 53884
rect 35076 53828 35080 53884
rect 35016 53824 35080 53828
rect 35096 53884 35160 53888
rect 35096 53828 35100 53884
rect 35100 53828 35156 53884
rect 35156 53828 35160 53884
rect 35096 53824 35160 53828
rect 35176 53884 35240 53888
rect 35176 53828 35180 53884
rect 35180 53828 35236 53884
rect 35236 53828 35240 53884
rect 35176 53824 35240 53828
rect 65656 53884 65720 53888
rect 65656 53828 65660 53884
rect 65660 53828 65716 53884
rect 65716 53828 65720 53884
rect 65656 53824 65720 53828
rect 65736 53884 65800 53888
rect 65736 53828 65740 53884
rect 65740 53828 65796 53884
rect 65796 53828 65800 53884
rect 65736 53824 65800 53828
rect 65816 53884 65880 53888
rect 65816 53828 65820 53884
rect 65820 53828 65876 53884
rect 65876 53828 65880 53884
rect 65816 53824 65880 53828
rect 65896 53884 65960 53888
rect 65896 53828 65900 53884
rect 65900 53828 65956 53884
rect 65956 53828 65960 53884
rect 65896 53824 65960 53828
rect 19576 53340 19640 53344
rect 19576 53284 19580 53340
rect 19580 53284 19636 53340
rect 19636 53284 19640 53340
rect 19576 53280 19640 53284
rect 19656 53340 19720 53344
rect 19656 53284 19660 53340
rect 19660 53284 19716 53340
rect 19716 53284 19720 53340
rect 19656 53280 19720 53284
rect 19736 53340 19800 53344
rect 19736 53284 19740 53340
rect 19740 53284 19796 53340
rect 19796 53284 19800 53340
rect 19736 53280 19800 53284
rect 19816 53340 19880 53344
rect 19816 53284 19820 53340
rect 19820 53284 19876 53340
rect 19876 53284 19880 53340
rect 19816 53280 19880 53284
rect 50296 53340 50360 53344
rect 50296 53284 50300 53340
rect 50300 53284 50356 53340
rect 50356 53284 50360 53340
rect 50296 53280 50360 53284
rect 50376 53340 50440 53344
rect 50376 53284 50380 53340
rect 50380 53284 50436 53340
rect 50436 53284 50440 53340
rect 50376 53280 50440 53284
rect 50456 53340 50520 53344
rect 50456 53284 50460 53340
rect 50460 53284 50516 53340
rect 50516 53284 50520 53340
rect 50456 53280 50520 53284
rect 50536 53340 50600 53344
rect 50536 53284 50540 53340
rect 50540 53284 50596 53340
rect 50596 53284 50600 53340
rect 50536 53280 50600 53284
rect 4216 52796 4280 52800
rect 4216 52740 4220 52796
rect 4220 52740 4276 52796
rect 4276 52740 4280 52796
rect 4216 52736 4280 52740
rect 4296 52796 4360 52800
rect 4296 52740 4300 52796
rect 4300 52740 4356 52796
rect 4356 52740 4360 52796
rect 4296 52736 4360 52740
rect 4376 52796 4440 52800
rect 4376 52740 4380 52796
rect 4380 52740 4436 52796
rect 4436 52740 4440 52796
rect 4376 52736 4440 52740
rect 4456 52796 4520 52800
rect 4456 52740 4460 52796
rect 4460 52740 4516 52796
rect 4516 52740 4520 52796
rect 4456 52736 4520 52740
rect 34936 52796 35000 52800
rect 34936 52740 34940 52796
rect 34940 52740 34996 52796
rect 34996 52740 35000 52796
rect 34936 52736 35000 52740
rect 35016 52796 35080 52800
rect 35016 52740 35020 52796
rect 35020 52740 35076 52796
rect 35076 52740 35080 52796
rect 35016 52736 35080 52740
rect 35096 52796 35160 52800
rect 35096 52740 35100 52796
rect 35100 52740 35156 52796
rect 35156 52740 35160 52796
rect 35096 52736 35160 52740
rect 35176 52796 35240 52800
rect 35176 52740 35180 52796
rect 35180 52740 35236 52796
rect 35236 52740 35240 52796
rect 35176 52736 35240 52740
rect 65656 52796 65720 52800
rect 65656 52740 65660 52796
rect 65660 52740 65716 52796
rect 65716 52740 65720 52796
rect 65656 52736 65720 52740
rect 65736 52796 65800 52800
rect 65736 52740 65740 52796
rect 65740 52740 65796 52796
rect 65796 52740 65800 52796
rect 65736 52736 65800 52740
rect 65816 52796 65880 52800
rect 65816 52740 65820 52796
rect 65820 52740 65876 52796
rect 65876 52740 65880 52796
rect 65816 52736 65880 52740
rect 65896 52796 65960 52800
rect 65896 52740 65900 52796
rect 65900 52740 65956 52796
rect 65956 52740 65960 52796
rect 65896 52736 65960 52740
rect 19576 52252 19640 52256
rect 19576 52196 19580 52252
rect 19580 52196 19636 52252
rect 19636 52196 19640 52252
rect 19576 52192 19640 52196
rect 19656 52252 19720 52256
rect 19656 52196 19660 52252
rect 19660 52196 19716 52252
rect 19716 52196 19720 52252
rect 19656 52192 19720 52196
rect 19736 52252 19800 52256
rect 19736 52196 19740 52252
rect 19740 52196 19796 52252
rect 19796 52196 19800 52252
rect 19736 52192 19800 52196
rect 19816 52252 19880 52256
rect 19816 52196 19820 52252
rect 19820 52196 19876 52252
rect 19876 52196 19880 52252
rect 19816 52192 19880 52196
rect 50296 52252 50360 52256
rect 50296 52196 50300 52252
rect 50300 52196 50356 52252
rect 50356 52196 50360 52252
rect 50296 52192 50360 52196
rect 50376 52252 50440 52256
rect 50376 52196 50380 52252
rect 50380 52196 50436 52252
rect 50436 52196 50440 52252
rect 50376 52192 50440 52196
rect 50456 52252 50520 52256
rect 50456 52196 50460 52252
rect 50460 52196 50516 52252
rect 50516 52196 50520 52252
rect 50456 52192 50520 52196
rect 50536 52252 50600 52256
rect 50536 52196 50540 52252
rect 50540 52196 50596 52252
rect 50596 52196 50600 52252
rect 50536 52192 50600 52196
rect 4216 51708 4280 51712
rect 4216 51652 4220 51708
rect 4220 51652 4276 51708
rect 4276 51652 4280 51708
rect 4216 51648 4280 51652
rect 4296 51708 4360 51712
rect 4296 51652 4300 51708
rect 4300 51652 4356 51708
rect 4356 51652 4360 51708
rect 4296 51648 4360 51652
rect 4376 51708 4440 51712
rect 4376 51652 4380 51708
rect 4380 51652 4436 51708
rect 4436 51652 4440 51708
rect 4376 51648 4440 51652
rect 4456 51708 4520 51712
rect 4456 51652 4460 51708
rect 4460 51652 4516 51708
rect 4516 51652 4520 51708
rect 4456 51648 4520 51652
rect 34936 51708 35000 51712
rect 34936 51652 34940 51708
rect 34940 51652 34996 51708
rect 34996 51652 35000 51708
rect 34936 51648 35000 51652
rect 35016 51708 35080 51712
rect 35016 51652 35020 51708
rect 35020 51652 35076 51708
rect 35076 51652 35080 51708
rect 35016 51648 35080 51652
rect 35096 51708 35160 51712
rect 35096 51652 35100 51708
rect 35100 51652 35156 51708
rect 35156 51652 35160 51708
rect 35096 51648 35160 51652
rect 35176 51708 35240 51712
rect 35176 51652 35180 51708
rect 35180 51652 35236 51708
rect 35236 51652 35240 51708
rect 35176 51648 35240 51652
rect 65656 51708 65720 51712
rect 65656 51652 65660 51708
rect 65660 51652 65716 51708
rect 65716 51652 65720 51708
rect 65656 51648 65720 51652
rect 65736 51708 65800 51712
rect 65736 51652 65740 51708
rect 65740 51652 65796 51708
rect 65796 51652 65800 51708
rect 65736 51648 65800 51652
rect 65816 51708 65880 51712
rect 65816 51652 65820 51708
rect 65820 51652 65876 51708
rect 65876 51652 65880 51708
rect 65816 51648 65880 51652
rect 65896 51708 65960 51712
rect 65896 51652 65900 51708
rect 65900 51652 65956 51708
rect 65956 51652 65960 51708
rect 65896 51648 65960 51652
rect 19576 51164 19640 51168
rect 19576 51108 19580 51164
rect 19580 51108 19636 51164
rect 19636 51108 19640 51164
rect 19576 51104 19640 51108
rect 19656 51164 19720 51168
rect 19656 51108 19660 51164
rect 19660 51108 19716 51164
rect 19716 51108 19720 51164
rect 19656 51104 19720 51108
rect 19736 51164 19800 51168
rect 19736 51108 19740 51164
rect 19740 51108 19796 51164
rect 19796 51108 19800 51164
rect 19736 51104 19800 51108
rect 19816 51164 19880 51168
rect 19816 51108 19820 51164
rect 19820 51108 19876 51164
rect 19876 51108 19880 51164
rect 19816 51104 19880 51108
rect 50296 51164 50360 51168
rect 50296 51108 50300 51164
rect 50300 51108 50356 51164
rect 50356 51108 50360 51164
rect 50296 51104 50360 51108
rect 50376 51164 50440 51168
rect 50376 51108 50380 51164
rect 50380 51108 50436 51164
rect 50436 51108 50440 51164
rect 50376 51104 50440 51108
rect 50456 51164 50520 51168
rect 50456 51108 50460 51164
rect 50460 51108 50516 51164
rect 50516 51108 50520 51164
rect 50456 51104 50520 51108
rect 50536 51164 50600 51168
rect 50536 51108 50540 51164
rect 50540 51108 50596 51164
rect 50596 51108 50600 51164
rect 50536 51104 50600 51108
rect 4216 50620 4280 50624
rect 4216 50564 4220 50620
rect 4220 50564 4276 50620
rect 4276 50564 4280 50620
rect 4216 50560 4280 50564
rect 4296 50620 4360 50624
rect 4296 50564 4300 50620
rect 4300 50564 4356 50620
rect 4356 50564 4360 50620
rect 4296 50560 4360 50564
rect 4376 50620 4440 50624
rect 4376 50564 4380 50620
rect 4380 50564 4436 50620
rect 4436 50564 4440 50620
rect 4376 50560 4440 50564
rect 4456 50620 4520 50624
rect 4456 50564 4460 50620
rect 4460 50564 4516 50620
rect 4516 50564 4520 50620
rect 4456 50560 4520 50564
rect 34936 50620 35000 50624
rect 34936 50564 34940 50620
rect 34940 50564 34996 50620
rect 34996 50564 35000 50620
rect 34936 50560 35000 50564
rect 35016 50620 35080 50624
rect 35016 50564 35020 50620
rect 35020 50564 35076 50620
rect 35076 50564 35080 50620
rect 35016 50560 35080 50564
rect 35096 50620 35160 50624
rect 35096 50564 35100 50620
rect 35100 50564 35156 50620
rect 35156 50564 35160 50620
rect 35096 50560 35160 50564
rect 35176 50620 35240 50624
rect 35176 50564 35180 50620
rect 35180 50564 35236 50620
rect 35236 50564 35240 50620
rect 35176 50560 35240 50564
rect 65656 50620 65720 50624
rect 65656 50564 65660 50620
rect 65660 50564 65716 50620
rect 65716 50564 65720 50620
rect 65656 50560 65720 50564
rect 65736 50620 65800 50624
rect 65736 50564 65740 50620
rect 65740 50564 65796 50620
rect 65796 50564 65800 50620
rect 65736 50560 65800 50564
rect 65816 50620 65880 50624
rect 65816 50564 65820 50620
rect 65820 50564 65876 50620
rect 65876 50564 65880 50620
rect 65816 50560 65880 50564
rect 65896 50620 65960 50624
rect 65896 50564 65900 50620
rect 65900 50564 65956 50620
rect 65956 50564 65960 50620
rect 65896 50560 65960 50564
rect 19576 50076 19640 50080
rect 19576 50020 19580 50076
rect 19580 50020 19636 50076
rect 19636 50020 19640 50076
rect 19576 50016 19640 50020
rect 19656 50076 19720 50080
rect 19656 50020 19660 50076
rect 19660 50020 19716 50076
rect 19716 50020 19720 50076
rect 19656 50016 19720 50020
rect 19736 50076 19800 50080
rect 19736 50020 19740 50076
rect 19740 50020 19796 50076
rect 19796 50020 19800 50076
rect 19736 50016 19800 50020
rect 19816 50076 19880 50080
rect 19816 50020 19820 50076
rect 19820 50020 19876 50076
rect 19876 50020 19880 50076
rect 19816 50016 19880 50020
rect 50296 50076 50360 50080
rect 50296 50020 50300 50076
rect 50300 50020 50356 50076
rect 50356 50020 50360 50076
rect 50296 50016 50360 50020
rect 50376 50076 50440 50080
rect 50376 50020 50380 50076
rect 50380 50020 50436 50076
rect 50436 50020 50440 50076
rect 50376 50016 50440 50020
rect 50456 50076 50520 50080
rect 50456 50020 50460 50076
rect 50460 50020 50516 50076
rect 50516 50020 50520 50076
rect 50456 50016 50520 50020
rect 50536 50076 50600 50080
rect 50536 50020 50540 50076
rect 50540 50020 50596 50076
rect 50596 50020 50600 50076
rect 50536 50016 50600 50020
rect 4216 49532 4280 49536
rect 4216 49476 4220 49532
rect 4220 49476 4276 49532
rect 4276 49476 4280 49532
rect 4216 49472 4280 49476
rect 4296 49532 4360 49536
rect 4296 49476 4300 49532
rect 4300 49476 4356 49532
rect 4356 49476 4360 49532
rect 4296 49472 4360 49476
rect 4376 49532 4440 49536
rect 4376 49476 4380 49532
rect 4380 49476 4436 49532
rect 4436 49476 4440 49532
rect 4376 49472 4440 49476
rect 4456 49532 4520 49536
rect 4456 49476 4460 49532
rect 4460 49476 4516 49532
rect 4516 49476 4520 49532
rect 4456 49472 4520 49476
rect 34936 49532 35000 49536
rect 34936 49476 34940 49532
rect 34940 49476 34996 49532
rect 34996 49476 35000 49532
rect 34936 49472 35000 49476
rect 35016 49532 35080 49536
rect 35016 49476 35020 49532
rect 35020 49476 35076 49532
rect 35076 49476 35080 49532
rect 35016 49472 35080 49476
rect 35096 49532 35160 49536
rect 35096 49476 35100 49532
rect 35100 49476 35156 49532
rect 35156 49476 35160 49532
rect 35096 49472 35160 49476
rect 35176 49532 35240 49536
rect 35176 49476 35180 49532
rect 35180 49476 35236 49532
rect 35236 49476 35240 49532
rect 35176 49472 35240 49476
rect 65656 49532 65720 49536
rect 65656 49476 65660 49532
rect 65660 49476 65716 49532
rect 65716 49476 65720 49532
rect 65656 49472 65720 49476
rect 65736 49532 65800 49536
rect 65736 49476 65740 49532
rect 65740 49476 65796 49532
rect 65796 49476 65800 49532
rect 65736 49472 65800 49476
rect 65816 49532 65880 49536
rect 65816 49476 65820 49532
rect 65820 49476 65876 49532
rect 65876 49476 65880 49532
rect 65816 49472 65880 49476
rect 65896 49532 65960 49536
rect 65896 49476 65900 49532
rect 65900 49476 65956 49532
rect 65956 49476 65960 49532
rect 65896 49472 65960 49476
rect 19576 48988 19640 48992
rect 19576 48932 19580 48988
rect 19580 48932 19636 48988
rect 19636 48932 19640 48988
rect 19576 48928 19640 48932
rect 19656 48988 19720 48992
rect 19656 48932 19660 48988
rect 19660 48932 19716 48988
rect 19716 48932 19720 48988
rect 19656 48928 19720 48932
rect 19736 48988 19800 48992
rect 19736 48932 19740 48988
rect 19740 48932 19796 48988
rect 19796 48932 19800 48988
rect 19736 48928 19800 48932
rect 19816 48988 19880 48992
rect 19816 48932 19820 48988
rect 19820 48932 19876 48988
rect 19876 48932 19880 48988
rect 19816 48928 19880 48932
rect 50296 48988 50360 48992
rect 50296 48932 50300 48988
rect 50300 48932 50356 48988
rect 50356 48932 50360 48988
rect 50296 48928 50360 48932
rect 50376 48988 50440 48992
rect 50376 48932 50380 48988
rect 50380 48932 50436 48988
rect 50436 48932 50440 48988
rect 50376 48928 50440 48932
rect 50456 48988 50520 48992
rect 50456 48932 50460 48988
rect 50460 48932 50516 48988
rect 50516 48932 50520 48988
rect 50456 48928 50520 48932
rect 50536 48988 50600 48992
rect 50536 48932 50540 48988
rect 50540 48932 50596 48988
rect 50596 48932 50600 48988
rect 50536 48928 50600 48932
rect 4216 48444 4280 48448
rect 4216 48388 4220 48444
rect 4220 48388 4276 48444
rect 4276 48388 4280 48444
rect 4216 48384 4280 48388
rect 4296 48444 4360 48448
rect 4296 48388 4300 48444
rect 4300 48388 4356 48444
rect 4356 48388 4360 48444
rect 4296 48384 4360 48388
rect 4376 48444 4440 48448
rect 4376 48388 4380 48444
rect 4380 48388 4436 48444
rect 4436 48388 4440 48444
rect 4376 48384 4440 48388
rect 4456 48444 4520 48448
rect 4456 48388 4460 48444
rect 4460 48388 4516 48444
rect 4516 48388 4520 48444
rect 4456 48384 4520 48388
rect 34936 48444 35000 48448
rect 34936 48388 34940 48444
rect 34940 48388 34996 48444
rect 34996 48388 35000 48444
rect 34936 48384 35000 48388
rect 35016 48444 35080 48448
rect 35016 48388 35020 48444
rect 35020 48388 35076 48444
rect 35076 48388 35080 48444
rect 35016 48384 35080 48388
rect 35096 48444 35160 48448
rect 35096 48388 35100 48444
rect 35100 48388 35156 48444
rect 35156 48388 35160 48444
rect 35096 48384 35160 48388
rect 35176 48444 35240 48448
rect 35176 48388 35180 48444
rect 35180 48388 35236 48444
rect 35236 48388 35240 48444
rect 35176 48384 35240 48388
rect 65656 48444 65720 48448
rect 65656 48388 65660 48444
rect 65660 48388 65716 48444
rect 65716 48388 65720 48444
rect 65656 48384 65720 48388
rect 65736 48444 65800 48448
rect 65736 48388 65740 48444
rect 65740 48388 65796 48444
rect 65796 48388 65800 48444
rect 65736 48384 65800 48388
rect 65816 48444 65880 48448
rect 65816 48388 65820 48444
rect 65820 48388 65876 48444
rect 65876 48388 65880 48444
rect 65816 48384 65880 48388
rect 65896 48444 65960 48448
rect 65896 48388 65900 48444
rect 65900 48388 65956 48444
rect 65956 48388 65960 48444
rect 65896 48384 65960 48388
rect 19576 47900 19640 47904
rect 19576 47844 19580 47900
rect 19580 47844 19636 47900
rect 19636 47844 19640 47900
rect 19576 47840 19640 47844
rect 19656 47900 19720 47904
rect 19656 47844 19660 47900
rect 19660 47844 19716 47900
rect 19716 47844 19720 47900
rect 19656 47840 19720 47844
rect 19736 47900 19800 47904
rect 19736 47844 19740 47900
rect 19740 47844 19796 47900
rect 19796 47844 19800 47900
rect 19736 47840 19800 47844
rect 19816 47900 19880 47904
rect 19816 47844 19820 47900
rect 19820 47844 19876 47900
rect 19876 47844 19880 47900
rect 19816 47840 19880 47844
rect 50296 47900 50360 47904
rect 50296 47844 50300 47900
rect 50300 47844 50356 47900
rect 50356 47844 50360 47900
rect 50296 47840 50360 47844
rect 50376 47900 50440 47904
rect 50376 47844 50380 47900
rect 50380 47844 50436 47900
rect 50436 47844 50440 47900
rect 50376 47840 50440 47844
rect 50456 47900 50520 47904
rect 50456 47844 50460 47900
rect 50460 47844 50516 47900
rect 50516 47844 50520 47900
rect 50456 47840 50520 47844
rect 50536 47900 50600 47904
rect 50536 47844 50540 47900
rect 50540 47844 50596 47900
rect 50596 47844 50600 47900
rect 50536 47840 50600 47844
rect 4216 47356 4280 47360
rect 4216 47300 4220 47356
rect 4220 47300 4276 47356
rect 4276 47300 4280 47356
rect 4216 47296 4280 47300
rect 4296 47356 4360 47360
rect 4296 47300 4300 47356
rect 4300 47300 4356 47356
rect 4356 47300 4360 47356
rect 4296 47296 4360 47300
rect 4376 47356 4440 47360
rect 4376 47300 4380 47356
rect 4380 47300 4436 47356
rect 4436 47300 4440 47356
rect 4376 47296 4440 47300
rect 4456 47356 4520 47360
rect 4456 47300 4460 47356
rect 4460 47300 4516 47356
rect 4516 47300 4520 47356
rect 4456 47296 4520 47300
rect 34936 47356 35000 47360
rect 34936 47300 34940 47356
rect 34940 47300 34996 47356
rect 34996 47300 35000 47356
rect 34936 47296 35000 47300
rect 35016 47356 35080 47360
rect 35016 47300 35020 47356
rect 35020 47300 35076 47356
rect 35076 47300 35080 47356
rect 35016 47296 35080 47300
rect 35096 47356 35160 47360
rect 35096 47300 35100 47356
rect 35100 47300 35156 47356
rect 35156 47300 35160 47356
rect 35096 47296 35160 47300
rect 35176 47356 35240 47360
rect 35176 47300 35180 47356
rect 35180 47300 35236 47356
rect 35236 47300 35240 47356
rect 35176 47296 35240 47300
rect 65656 47356 65720 47360
rect 65656 47300 65660 47356
rect 65660 47300 65716 47356
rect 65716 47300 65720 47356
rect 65656 47296 65720 47300
rect 65736 47356 65800 47360
rect 65736 47300 65740 47356
rect 65740 47300 65796 47356
rect 65796 47300 65800 47356
rect 65736 47296 65800 47300
rect 65816 47356 65880 47360
rect 65816 47300 65820 47356
rect 65820 47300 65876 47356
rect 65876 47300 65880 47356
rect 65816 47296 65880 47300
rect 65896 47356 65960 47360
rect 65896 47300 65900 47356
rect 65900 47300 65956 47356
rect 65956 47300 65960 47356
rect 65896 47296 65960 47300
rect 19576 46812 19640 46816
rect 19576 46756 19580 46812
rect 19580 46756 19636 46812
rect 19636 46756 19640 46812
rect 19576 46752 19640 46756
rect 19656 46812 19720 46816
rect 19656 46756 19660 46812
rect 19660 46756 19716 46812
rect 19716 46756 19720 46812
rect 19656 46752 19720 46756
rect 19736 46812 19800 46816
rect 19736 46756 19740 46812
rect 19740 46756 19796 46812
rect 19796 46756 19800 46812
rect 19736 46752 19800 46756
rect 19816 46812 19880 46816
rect 19816 46756 19820 46812
rect 19820 46756 19876 46812
rect 19876 46756 19880 46812
rect 19816 46752 19880 46756
rect 50296 46812 50360 46816
rect 50296 46756 50300 46812
rect 50300 46756 50356 46812
rect 50356 46756 50360 46812
rect 50296 46752 50360 46756
rect 50376 46812 50440 46816
rect 50376 46756 50380 46812
rect 50380 46756 50436 46812
rect 50436 46756 50440 46812
rect 50376 46752 50440 46756
rect 50456 46812 50520 46816
rect 50456 46756 50460 46812
rect 50460 46756 50516 46812
rect 50516 46756 50520 46812
rect 50456 46752 50520 46756
rect 50536 46812 50600 46816
rect 50536 46756 50540 46812
rect 50540 46756 50596 46812
rect 50596 46756 50600 46812
rect 50536 46752 50600 46756
rect 4216 46268 4280 46272
rect 4216 46212 4220 46268
rect 4220 46212 4276 46268
rect 4276 46212 4280 46268
rect 4216 46208 4280 46212
rect 4296 46268 4360 46272
rect 4296 46212 4300 46268
rect 4300 46212 4356 46268
rect 4356 46212 4360 46268
rect 4296 46208 4360 46212
rect 4376 46268 4440 46272
rect 4376 46212 4380 46268
rect 4380 46212 4436 46268
rect 4436 46212 4440 46268
rect 4376 46208 4440 46212
rect 4456 46268 4520 46272
rect 4456 46212 4460 46268
rect 4460 46212 4516 46268
rect 4516 46212 4520 46268
rect 4456 46208 4520 46212
rect 34936 46268 35000 46272
rect 34936 46212 34940 46268
rect 34940 46212 34996 46268
rect 34996 46212 35000 46268
rect 34936 46208 35000 46212
rect 35016 46268 35080 46272
rect 35016 46212 35020 46268
rect 35020 46212 35076 46268
rect 35076 46212 35080 46268
rect 35016 46208 35080 46212
rect 35096 46268 35160 46272
rect 35096 46212 35100 46268
rect 35100 46212 35156 46268
rect 35156 46212 35160 46268
rect 35096 46208 35160 46212
rect 35176 46268 35240 46272
rect 35176 46212 35180 46268
rect 35180 46212 35236 46268
rect 35236 46212 35240 46268
rect 35176 46208 35240 46212
rect 65656 46268 65720 46272
rect 65656 46212 65660 46268
rect 65660 46212 65716 46268
rect 65716 46212 65720 46268
rect 65656 46208 65720 46212
rect 65736 46268 65800 46272
rect 65736 46212 65740 46268
rect 65740 46212 65796 46268
rect 65796 46212 65800 46268
rect 65736 46208 65800 46212
rect 65816 46268 65880 46272
rect 65816 46212 65820 46268
rect 65820 46212 65876 46268
rect 65876 46212 65880 46268
rect 65816 46208 65880 46212
rect 65896 46268 65960 46272
rect 65896 46212 65900 46268
rect 65900 46212 65956 46268
rect 65956 46212 65960 46268
rect 65896 46208 65960 46212
rect 19576 45724 19640 45728
rect 19576 45668 19580 45724
rect 19580 45668 19636 45724
rect 19636 45668 19640 45724
rect 19576 45664 19640 45668
rect 19656 45724 19720 45728
rect 19656 45668 19660 45724
rect 19660 45668 19716 45724
rect 19716 45668 19720 45724
rect 19656 45664 19720 45668
rect 19736 45724 19800 45728
rect 19736 45668 19740 45724
rect 19740 45668 19796 45724
rect 19796 45668 19800 45724
rect 19736 45664 19800 45668
rect 19816 45724 19880 45728
rect 19816 45668 19820 45724
rect 19820 45668 19876 45724
rect 19876 45668 19880 45724
rect 19816 45664 19880 45668
rect 50296 45724 50360 45728
rect 50296 45668 50300 45724
rect 50300 45668 50356 45724
rect 50356 45668 50360 45724
rect 50296 45664 50360 45668
rect 50376 45724 50440 45728
rect 50376 45668 50380 45724
rect 50380 45668 50436 45724
rect 50436 45668 50440 45724
rect 50376 45664 50440 45668
rect 50456 45724 50520 45728
rect 50456 45668 50460 45724
rect 50460 45668 50516 45724
rect 50516 45668 50520 45724
rect 50456 45664 50520 45668
rect 50536 45724 50600 45728
rect 50536 45668 50540 45724
rect 50540 45668 50596 45724
rect 50596 45668 50600 45724
rect 50536 45664 50600 45668
rect 4216 45180 4280 45184
rect 4216 45124 4220 45180
rect 4220 45124 4276 45180
rect 4276 45124 4280 45180
rect 4216 45120 4280 45124
rect 4296 45180 4360 45184
rect 4296 45124 4300 45180
rect 4300 45124 4356 45180
rect 4356 45124 4360 45180
rect 4296 45120 4360 45124
rect 4376 45180 4440 45184
rect 4376 45124 4380 45180
rect 4380 45124 4436 45180
rect 4436 45124 4440 45180
rect 4376 45120 4440 45124
rect 4456 45180 4520 45184
rect 4456 45124 4460 45180
rect 4460 45124 4516 45180
rect 4516 45124 4520 45180
rect 4456 45120 4520 45124
rect 34936 45180 35000 45184
rect 34936 45124 34940 45180
rect 34940 45124 34996 45180
rect 34996 45124 35000 45180
rect 34936 45120 35000 45124
rect 35016 45180 35080 45184
rect 35016 45124 35020 45180
rect 35020 45124 35076 45180
rect 35076 45124 35080 45180
rect 35016 45120 35080 45124
rect 35096 45180 35160 45184
rect 35096 45124 35100 45180
rect 35100 45124 35156 45180
rect 35156 45124 35160 45180
rect 35096 45120 35160 45124
rect 35176 45180 35240 45184
rect 35176 45124 35180 45180
rect 35180 45124 35236 45180
rect 35236 45124 35240 45180
rect 35176 45120 35240 45124
rect 65656 45180 65720 45184
rect 65656 45124 65660 45180
rect 65660 45124 65716 45180
rect 65716 45124 65720 45180
rect 65656 45120 65720 45124
rect 65736 45180 65800 45184
rect 65736 45124 65740 45180
rect 65740 45124 65796 45180
rect 65796 45124 65800 45180
rect 65736 45120 65800 45124
rect 65816 45180 65880 45184
rect 65816 45124 65820 45180
rect 65820 45124 65876 45180
rect 65876 45124 65880 45180
rect 65816 45120 65880 45124
rect 65896 45180 65960 45184
rect 65896 45124 65900 45180
rect 65900 45124 65956 45180
rect 65956 45124 65960 45180
rect 65896 45120 65960 45124
rect 19576 44636 19640 44640
rect 19576 44580 19580 44636
rect 19580 44580 19636 44636
rect 19636 44580 19640 44636
rect 19576 44576 19640 44580
rect 19656 44636 19720 44640
rect 19656 44580 19660 44636
rect 19660 44580 19716 44636
rect 19716 44580 19720 44636
rect 19656 44576 19720 44580
rect 19736 44636 19800 44640
rect 19736 44580 19740 44636
rect 19740 44580 19796 44636
rect 19796 44580 19800 44636
rect 19736 44576 19800 44580
rect 19816 44636 19880 44640
rect 19816 44580 19820 44636
rect 19820 44580 19876 44636
rect 19876 44580 19880 44636
rect 19816 44576 19880 44580
rect 50296 44636 50360 44640
rect 50296 44580 50300 44636
rect 50300 44580 50356 44636
rect 50356 44580 50360 44636
rect 50296 44576 50360 44580
rect 50376 44636 50440 44640
rect 50376 44580 50380 44636
rect 50380 44580 50436 44636
rect 50436 44580 50440 44636
rect 50376 44576 50440 44580
rect 50456 44636 50520 44640
rect 50456 44580 50460 44636
rect 50460 44580 50516 44636
rect 50516 44580 50520 44636
rect 50456 44576 50520 44580
rect 50536 44636 50600 44640
rect 50536 44580 50540 44636
rect 50540 44580 50596 44636
rect 50596 44580 50600 44636
rect 50536 44576 50600 44580
rect 4216 44092 4280 44096
rect 4216 44036 4220 44092
rect 4220 44036 4276 44092
rect 4276 44036 4280 44092
rect 4216 44032 4280 44036
rect 4296 44092 4360 44096
rect 4296 44036 4300 44092
rect 4300 44036 4356 44092
rect 4356 44036 4360 44092
rect 4296 44032 4360 44036
rect 4376 44092 4440 44096
rect 4376 44036 4380 44092
rect 4380 44036 4436 44092
rect 4436 44036 4440 44092
rect 4376 44032 4440 44036
rect 4456 44092 4520 44096
rect 4456 44036 4460 44092
rect 4460 44036 4516 44092
rect 4516 44036 4520 44092
rect 4456 44032 4520 44036
rect 34936 44092 35000 44096
rect 34936 44036 34940 44092
rect 34940 44036 34996 44092
rect 34996 44036 35000 44092
rect 34936 44032 35000 44036
rect 35016 44092 35080 44096
rect 35016 44036 35020 44092
rect 35020 44036 35076 44092
rect 35076 44036 35080 44092
rect 35016 44032 35080 44036
rect 35096 44092 35160 44096
rect 35096 44036 35100 44092
rect 35100 44036 35156 44092
rect 35156 44036 35160 44092
rect 35096 44032 35160 44036
rect 35176 44092 35240 44096
rect 35176 44036 35180 44092
rect 35180 44036 35236 44092
rect 35236 44036 35240 44092
rect 35176 44032 35240 44036
rect 65656 44092 65720 44096
rect 65656 44036 65660 44092
rect 65660 44036 65716 44092
rect 65716 44036 65720 44092
rect 65656 44032 65720 44036
rect 65736 44092 65800 44096
rect 65736 44036 65740 44092
rect 65740 44036 65796 44092
rect 65796 44036 65800 44092
rect 65736 44032 65800 44036
rect 65816 44092 65880 44096
rect 65816 44036 65820 44092
rect 65820 44036 65876 44092
rect 65876 44036 65880 44092
rect 65816 44032 65880 44036
rect 65896 44092 65960 44096
rect 65896 44036 65900 44092
rect 65900 44036 65956 44092
rect 65956 44036 65960 44092
rect 65896 44032 65960 44036
rect 19576 43548 19640 43552
rect 19576 43492 19580 43548
rect 19580 43492 19636 43548
rect 19636 43492 19640 43548
rect 19576 43488 19640 43492
rect 19656 43548 19720 43552
rect 19656 43492 19660 43548
rect 19660 43492 19716 43548
rect 19716 43492 19720 43548
rect 19656 43488 19720 43492
rect 19736 43548 19800 43552
rect 19736 43492 19740 43548
rect 19740 43492 19796 43548
rect 19796 43492 19800 43548
rect 19736 43488 19800 43492
rect 19816 43548 19880 43552
rect 19816 43492 19820 43548
rect 19820 43492 19876 43548
rect 19876 43492 19880 43548
rect 19816 43488 19880 43492
rect 50296 43548 50360 43552
rect 50296 43492 50300 43548
rect 50300 43492 50356 43548
rect 50356 43492 50360 43548
rect 50296 43488 50360 43492
rect 50376 43548 50440 43552
rect 50376 43492 50380 43548
rect 50380 43492 50436 43548
rect 50436 43492 50440 43548
rect 50376 43488 50440 43492
rect 50456 43548 50520 43552
rect 50456 43492 50460 43548
rect 50460 43492 50516 43548
rect 50516 43492 50520 43548
rect 50456 43488 50520 43492
rect 50536 43548 50600 43552
rect 50536 43492 50540 43548
rect 50540 43492 50596 43548
rect 50596 43492 50600 43548
rect 50536 43488 50600 43492
rect 4216 43004 4280 43008
rect 4216 42948 4220 43004
rect 4220 42948 4276 43004
rect 4276 42948 4280 43004
rect 4216 42944 4280 42948
rect 4296 43004 4360 43008
rect 4296 42948 4300 43004
rect 4300 42948 4356 43004
rect 4356 42948 4360 43004
rect 4296 42944 4360 42948
rect 4376 43004 4440 43008
rect 4376 42948 4380 43004
rect 4380 42948 4436 43004
rect 4436 42948 4440 43004
rect 4376 42944 4440 42948
rect 4456 43004 4520 43008
rect 4456 42948 4460 43004
rect 4460 42948 4516 43004
rect 4516 42948 4520 43004
rect 4456 42944 4520 42948
rect 34936 43004 35000 43008
rect 34936 42948 34940 43004
rect 34940 42948 34996 43004
rect 34996 42948 35000 43004
rect 34936 42944 35000 42948
rect 35016 43004 35080 43008
rect 35016 42948 35020 43004
rect 35020 42948 35076 43004
rect 35076 42948 35080 43004
rect 35016 42944 35080 42948
rect 35096 43004 35160 43008
rect 35096 42948 35100 43004
rect 35100 42948 35156 43004
rect 35156 42948 35160 43004
rect 35096 42944 35160 42948
rect 35176 43004 35240 43008
rect 35176 42948 35180 43004
rect 35180 42948 35236 43004
rect 35236 42948 35240 43004
rect 35176 42944 35240 42948
rect 65656 43004 65720 43008
rect 65656 42948 65660 43004
rect 65660 42948 65716 43004
rect 65716 42948 65720 43004
rect 65656 42944 65720 42948
rect 65736 43004 65800 43008
rect 65736 42948 65740 43004
rect 65740 42948 65796 43004
rect 65796 42948 65800 43004
rect 65736 42944 65800 42948
rect 65816 43004 65880 43008
rect 65816 42948 65820 43004
rect 65820 42948 65876 43004
rect 65876 42948 65880 43004
rect 65816 42944 65880 42948
rect 65896 43004 65960 43008
rect 65896 42948 65900 43004
rect 65900 42948 65956 43004
rect 65956 42948 65960 43004
rect 65896 42944 65960 42948
rect 19576 42460 19640 42464
rect 19576 42404 19580 42460
rect 19580 42404 19636 42460
rect 19636 42404 19640 42460
rect 19576 42400 19640 42404
rect 19656 42460 19720 42464
rect 19656 42404 19660 42460
rect 19660 42404 19716 42460
rect 19716 42404 19720 42460
rect 19656 42400 19720 42404
rect 19736 42460 19800 42464
rect 19736 42404 19740 42460
rect 19740 42404 19796 42460
rect 19796 42404 19800 42460
rect 19736 42400 19800 42404
rect 19816 42460 19880 42464
rect 19816 42404 19820 42460
rect 19820 42404 19876 42460
rect 19876 42404 19880 42460
rect 19816 42400 19880 42404
rect 50296 42460 50360 42464
rect 50296 42404 50300 42460
rect 50300 42404 50356 42460
rect 50356 42404 50360 42460
rect 50296 42400 50360 42404
rect 50376 42460 50440 42464
rect 50376 42404 50380 42460
rect 50380 42404 50436 42460
rect 50436 42404 50440 42460
rect 50376 42400 50440 42404
rect 50456 42460 50520 42464
rect 50456 42404 50460 42460
rect 50460 42404 50516 42460
rect 50516 42404 50520 42460
rect 50456 42400 50520 42404
rect 50536 42460 50600 42464
rect 50536 42404 50540 42460
rect 50540 42404 50596 42460
rect 50596 42404 50600 42460
rect 50536 42400 50600 42404
rect 4216 41916 4280 41920
rect 4216 41860 4220 41916
rect 4220 41860 4276 41916
rect 4276 41860 4280 41916
rect 4216 41856 4280 41860
rect 4296 41916 4360 41920
rect 4296 41860 4300 41916
rect 4300 41860 4356 41916
rect 4356 41860 4360 41916
rect 4296 41856 4360 41860
rect 4376 41916 4440 41920
rect 4376 41860 4380 41916
rect 4380 41860 4436 41916
rect 4436 41860 4440 41916
rect 4376 41856 4440 41860
rect 4456 41916 4520 41920
rect 4456 41860 4460 41916
rect 4460 41860 4516 41916
rect 4516 41860 4520 41916
rect 4456 41856 4520 41860
rect 34936 41916 35000 41920
rect 34936 41860 34940 41916
rect 34940 41860 34996 41916
rect 34996 41860 35000 41916
rect 34936 41856 35000 41860
rect 35016 41916 35080 41920
rect 35016 41860 35020 41916
rect 35020 41860 35076 41916
rect 35076 41860 35080 41916
rect 35016 41856 35080 41860
rect 35096 41916 35160 41920
rect 35096 41860 35100 41916
rect 35100 41860 35156 41916
rect 35156 41860 35160 41916
rect 35096 41856 35160 41860
rect 35176 41916 35240 41920
rect 35176 41860 35180 41916
rect 35180 41860 35236 41916
rect 35236 41860 35240 41916
rect 35176 41856 35240 41860
rect 65656 41916 65720 41920
rect 65656 41860 65660 41916
rect 65660 41860 65716 41916
rect 65716 41860 65720 41916
rect 65656 41856 65720 41860
rect 65736 41916 65800 41920
rect 65736 41860 65740 41916
rect 65740 41860 65796 41916
rect 65796 41860 65800 41916
rect 65736 41856 65800 41860
rect 65816 41916 65880 41920
rect 65816 41860 65820 41916
rect 65820 41860 65876 41916
rect 65876 41860 65880 41916
rect 65816 41856 65880 41860
rect 65896 41916 65960 41920
rect 65896 41860 65900 41916
rect 65900 41860 65956 41916
rect 65956 41860 65960 41916
rect 65896 41856 65960 41860
rect 19576 41372 19640 41376
rect 19576 41316 19580 41372
rect 19580 41316 19636 41372
rect 19636 41316 19640 41372
rect 19576 41312 19640 41316
rect 19656 41372 19720 41376
rect 19656 41316 19660 41372
rect 19660 41316 19716 41372
rect 19716 41316 19720 41372
rect 19656 41312 19720 41316
rect 19736 41372 19800 41376
rect 19736 41316 19740 41372
rect 19740 41316 19796 41372
rect 19796 41316 19800 41372
rect 19736 41312 19800 41316
rect 19816 41372 19880 41376
rect 19816 41316 19820 41372
rect 19820 41316 19876 41372
rect 19876 41316 19880 41372
rect 19816 41312 19880 41316
rect 50296 41372 50360 41376
rect 50296 41316 50300 41372
rect 50300 41316 50356 41372
rect 50356 41316 50360 41372
rect 50296 41312 50360 41316
rect 50376 41372 50440 41376
rect 50376 41316 50380 41372
rect 50380 41316 50436 41372
rect 50436 41316 50440 41372
rect 50376 41312 50440 41316
rect 50456 41372 50520 41376
rect 50456 41316 50460 41372
rect 50460 41316 50516 41372
rect 50516 41316 50520 41372
rect 50456 41312 50520 41316
rect 50536 41372 50600 41376
rect 50536 41316 50540 41372
rect 50540 41316 50596 41372
rect 50596 41316 50600 41372
rect 50536 41312 50600 41316
rect 4216 40828 4280 40832
rect 4216 40772 4220 40828
rect 4220 40772 4276 40828
rect 4276 40772 4280 40828
rect 4216 40768 4280 40772
rect 4296 40828 4360 40832
rect 4296 40772 4300 40828
rect 4300 40772 4356 40828
rect 4356 40772 4360 40828
rect 4296 40768 4360 40772
rect 4376 40828 4440 40832
rect 4376 40772 4380 40828
rect 4380 40772 4436 40828
rect 4436 40772 4440 40828
rect 4376 40768 4440 40772
rect 4456 40828 4520 40832
rect 4456 40772 4460 40828
rect 4460 40772 4516 40828
rect 4516 40772 4520 40828
rect 4456 40768 4520 40772
rect 34936 40828 35000 40832
rect 34936 40772 34940 40828
rect 34940 40772 34996 40828
rect 34996 40772 35000 40828
rect 34936 40768 35000 40772
rect 35016 40828 35080 40832
rect 35016 40772 35020 40828
rect 35020 40772 35076 40828
rect 35076 40772 35080 40828
rect 35016 40768 35080 40772
rect 35096 40828 35160 40832
rect 35096 40772 35100 40828
rect 35100 40772 35156 40828
rect 35156 40772 35160 40828
rect 35096 40768 35160 40772
rect 35176 40828 35240 40832
rect 35176 40772 35180 40828
rect 35180 40772 35236 40828
rect 35236 40772 35240 40828
rect 35176 40768 35240 40772
rect 65656 40828 65720 40832
rect 65656 40772 65660 40828
rect 65660 40772 65716 40828
rect 65716 40772 65720 40828
rect 65656 40768 65720 40772
rect 65736 40828 65800 40832
rect 65736 40772 65740 40828
rect 65740 40772 65796 40828
rect 65796 40772 65800 40828
rect 65736 40768 65800 40772
rect 65816 40828 65880 40832
rect 65816 40772 65820 40828
rect 65820 40772 65876 40828
rect 65876 40772 65880 40828
rect 65816 40768 65880 40772
rect 65896 40828 65960 40832
rect 65896 40772 65900 40828
rect 65900 40772 65956 40828
rect 65956 40772 65960 40828
rect 65896 40768 65960 40772
rect 19576 40284 19640 40288
rect 19576 40228 19580 40284
rect 19580 40228 19636 40284
rect 19636 40228 19640 40284
rect 19576 40224 19640 40228
rect 19656 40284 19720 40288
rect 19656 40228 19660 40284
rect 19660 40228 19716 40284
rect 19716 40228 19720 40284
rect 19656 40224 19720 40228
rect 19736 40284 19800 40288
rect 19736 40228 19740 40284
rect 19740 40228 19796 40284
rect 19796 40228 19800 40284
rect 19736 40224 19800 40228
rect 19816 40284 19880 40288
rect 19816 40228 19820 40284
rect 19820 40228 19876 40284
rect 19876 40228 19880 40284
rect 19816 40224 19880 40228
rect 50296 40284 50360 40288
rect 50296 40228 50300 40284
rect 50300 40228 50356 40284
rect 50356 40228 50360 40284
rect 50296 40224 50360 40228
rect 50376 40284 50440 40288
rect 50376 40228 50380 40284
rect 50380 40228 50436 40284
rect 50436 40228 50440 40284
rect 50376 40224 50440 40228
rect 50456 40284 50520 40288
rect 50456 40228 50460 40284
rect 50460 40228 50516 40284
rect 50516 40228 50520 40284
rect 50456 40224 50520 40228
rect 50536 40284 50600 40288
rect 50536 40228 50540 40284
rect 50540 40228 50596 40284
rect 50596 40228 50600 40284
rect 50536 40224 50600 40228
rect 4216 39740 4280 39744
rect 4216 39684 4220 39740
rect 4220 39684 4276 39740
rect 4276 39684 4280 39740
rect 4216 39680 4280 39684
rect 4296 39740 4360 39744
rect 4296 39684 4300 39740
rect 4300 39684 4356 39740
rect 4356 39684 4360 39740
rect 4296 39680 4360 39684
rect 4376 39740 4440 39744
rect 4376 39684 4380 39740
rect 4380 39684 4436 39740
rect 4436 39684 4440 39740
rect 4376 39680 4440 39684
rect 4456 39740 4520 39744
rect 4456 39684 4460 39740
rect 4460 39684 4516 39740
rect 4516 39684 4520 39740
rect 4456 39680 4520 39684
rect 34936 39740 35000 39744
rect 34936 39684 34940 39740
rect 34940 39684 34996 39740
rect 34996 39684 35000 39740
rect 34936 39680 35000 39684
rect 35016 39740 35080 39744
rect 35016 39684 35020 39740
rect 35020 39684 35076 39740
rect 35076 39684 35080 39740
rect 35016 39680 35080 39684
rect 35096 39740 35160 39744
rect 35096 39684 35100 39740
rect 35100 39684 35156 39740
rect 35156 39684 35160 39740
rect 35096 39680 35160 39684
rect 35176 39740 35240 39744
rect 35176 39684 35180 39740
rect 35180 39684 35236 39740
rect 35236 39684 35240 39740
rect 35176 39680 35240 39684
rect 65656 39740 65720 39744
rect 65656 39684 65660 39740
rect 65660 39684 65716 39740
rect 65716 39684 65720 39740
rect 65656 39680 65720 39684
rect 65736 39740 65800 39744
rect 65736 39684 65740 39740
rect 65740 39684 65796 39740
rect 65796 39684 65800 39740
rect 65736 39680 65800 39684
rect 65816 39740 65880 39744
rect 65816 39684 65820 39740
rect 65820 39684 65876 39740
rect 65876 39684 65880 39740
rect 65816 39680 65880 39684
rect 65896 39740 65960 39744
rect 65896 39684 65900 39740
rect 65900 39684 65956 39740
rect 65956 39684 65960 39740
rect 65896 39680 65960 39684
rect 19576 39196 19640 39200
rect 19576 39140 19580 39196
rect 19580 39140 19636 39196
rect 19636 39140 19640 39196
rect 19576 39136 19640 39140
rect 19656 39196 19720 39200
rect 19656 39140 19660 39196
rect 19660 39140 19716 39196
rect 19716 39140 19720 39196
rect 19656 39136 19720 39140
rect 19736 39196 19800 39200
rect 19736 39140 19740 39196
rect 19740 39140 19796 39196
rect 19796 39140 19800 39196
rect 19736 39136 19800 39140
rect 19816 39196 19880 39200
rect 19816 39140 19820 39196
rect 19820 39140 19876 39196
rect 19876 39140 19880 39196
rect 19816 39136 19880 39140
rect 50296 39196 50360 39200
rect 50296 39140 50300 39196
rect 50300 39140 50356 39196
rect 50356 39140 50360 39196
rect 50296 39136 50360 39140
rect 50376 39196 50440 39200
rect 50376 39140 50380 39196
rect 50380 39140 50436 39196
rect 50436 39140 50440 39196
rect 50376 39136 50440 39140
rect 50456 39196 50520 39200
rect 50456 39140 50460 39196
rect 50460 39140 50516 39196
rect 50516 39140 50520 39196
rect 50456 39136 50520 39140
rect 50536 39196 50600 39200
rect 50536 39140 50540 39196
rect 50540 39140 50596 39196
rect 50596 39140 50600 39196
rect 50536 39136 50600 39140
rect 4216 38652 4280 38656
rect 4216 38596 4220 38652
rect 4220 38596 4276 38652
rect 4276 38596 4280 38652
rect 4216 38592 4280 38596
rect 4296 38652 4360 38656
rect 4296 38596 4300 38652
rect 4300 38596 4356 38652
rect 4356 38596 4360 38652
rect 4296 38592 4360 38596
rect 4376 38652 4440 38656
rect 4376 38596 4380 38652
rect 4380 38596 4436 38652
rect 4436 38596 4440 38652
rect 4376 38592 4440 38596
rect 4456 38652 4520 38656
rect 4456 38596 4460 38652
rect 4460 38596 4516 38652
rect 4516 38596 4520 38652
rect 4456 38592 4520 38596
rect 34936 38652 35000 38656
rect 34936 38596 34940 38652
rect 34940 38596 34996 38652
rect 34996 38596 35000 38652
rect 34936 38592 35000 38596
rect 35016 38652 35080 38656
rect 35016 38596 35020 38652
rect 35020 38596 35076 38652
rect 35076 38596 35080 38652
rect 35016 38592 35080 38596
rect 35096 38652 35160 38656
rect 35096 38596 35100 38652
rect 35100 38596 35156 38652
rect 35156 38596 35160 38652
rect 35096 38592 35160 38596
rect 35176 38652 35240 38656
rect 35176 38596 35180 38652
rect 35180 38596 35236 38652
rect 35236 38596 35240 38652
rect 35176 38592 35240 38596
rect 65656 38652 65720 38656
rect 65656 38596 65660 38652
rect 65660 38596 65716 38652
rect 65716 38596 65720 38652
rect 65656 38592 65720 38596
rect 65736 38652 65800 38656
rect 65736 38596 65740 38652
rect 65740 38596 65796 38652
rect 65796 38596 65800 38652
rect 65736 38592 65800 38596
rect 65816 38652 65880 38656
rect 65816 38596 65820 38652
rect 65820 38596 65876 38652
rect 65876 38596 65880 38652
rect 65816 38592 65880 38596
rect 65896 38652 65960 38656
rect 65896 38596 65900 38652
rect 65900 38596 65956 38652
rect 65956 38596 65960 38652
rect 65896 38592 65960 38596
rect 19576 38108 19640 38112
rect 19576 38052 19580 38108
rect 19580 38052 19636 38108
rect 19636 38052 19640 38108
rect 19576 38048 19640 38052
rect 19656 38108 19720 38112
rect 19656 38052 19660 38108
rect 19660 38052 19716 38108
rect 19716 38052 19720 38108
rect 19656 38048 19720 38052
rect 19736 38108 19800 38112
rect 19736 38052 19740 38108
rect 19740 38052 19796 38108
rect 19796 38052 19800 38108
rect 19736 38048 19800 38052
rect 19816 38108 19880 38112
rect 19816 38052 19820 38108
rect 19820 38052 19876 38108
rect 19876 38052 19880 38108
rect 19816 38048 19880 38052
rect 50296 38108 50360 38112
rect 50296 38052 50300 38108
rect 50300 38052 50356 38108
rect 50356 38052 50360 38108
rect 50296 38048 50360 38052
rect 50376 38108 50440 38112
rect 50376 38052 50380 38108
rect 50380 38052 50436 38108
rect 50436 38052 50440 38108
rect 50376 38048 50440 38052
rect 50456 38108 50520 38112
rect 50456 38052 50460 38108
rect 50460 38052 50516 38108
rect 50516 38052 50520 38108
rect 50456 38048 50520 38052
rect 50536 38108 50600 38112
rect 50536 38052 50540 38108
rect 50540 38052 50596 38108
rect 50596 38052 50600 38108
rect 50536 38048 50600 38052
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 34936 37564 35000 37568
rect 34936 37508 34940 37564
rect 34940 37508 34996 37564
rect 34996 37508 35000 37564
rect 34936 37504 35000 37508
rect 35016 37564 35080 37568
rect 35016 37508 35020 37564
rect 35020 37508 35076 37564
rect 35076 37508 35080 37564
rect 35016 37504 35080 37508
rect 35096 37564 35160 37568
rect 35096 37508 35100 37564
rect 35100 37508 35156 37564
rect 35156 37508 35160 37564
rect 35096 37504 35160 37508
rect 35176 37564 35240 37568
rect 35176 37508 35180 37564
rect 35180 37508 35236 37564
rect 35236 37508 35240 37564
rect 35176 37504 35240 37508
rect 65656 37564 65720 37568
rect 65656 37508 65660 37564
rect 65660 37508 65716 37564
rect 65716 37508 65720 37564
rect 65656 37504 65720 37508
rect 65736 37564 65800 37568
rect 65736 37508 65740 37564
rect 65740 37508 65796 37564
rect 65796 37508 65800 37564
rect 65736 37504 65800 37508
rect 65816 37564 65880 37568
rect 65816 37508 65820 37564
rect 65820 37508 65876 37564
rect 65876 37508 65880 37564
rect 65816 37504 65880 37508
rect 65896 37564 65960 37568
rect 65896 37508 65900 37564
rect 65900 37508 65956 37564
rect 65956 37508 65960 37564
rect 65896 37504 65960 37508
rect 19576 37020 19640 37024
rect 19576 36964 19580 37020
rect 19580 36964 19636 37020
rect 19636 36964 19640 37020
rect 19576 36960 19640 36964
rect 19656 37020 19720 37024
rect 19656 36964 19660 37020
rect 19660 36964 19716 37020
rect 19716 36964 19720 37020
rect 19656 36960 19720 36964
rect 19736 37020 19800 37024
rect 19736 36964 19740 37020
rect 19740 36964 19796 37020
rect 19796 36964 19800 37020
rect 19736 36960 19800 36964
rect 19816 37020 19880 37024
rect 19816 36964 19820 37020
rect 19820 36964 19876 37020
rect 19876 36964 19880 37020
rect 19816 36960 19880 36964
rect 50296 37020 50360 37024
rect 50296 36964 50300 37020
rect 50300 36964 50356 37020
rect 50356 36964 50360 37020
rect 50296 36960 50360 36964
rect 50376 37020 50440 37024
rect 50376 36964 50380 37020
rect 50380 36964 50436 37020
rect 50436 36964 50440 37020
rect 50376 36960 50440 36964
rect 50456 37020 50520 37024
rect 50456 36964 50460 37020
rect 50460 36964 50516 37020
rect 50516 36964 50520 37020
rect 50456 36960 50520 36964
rect 50536 37020 50600 37024
rect 50536 36964 50540 37020
rect 50540 36964 50596 37020
rect 50596 36964 50600 37020
rect 50536 36960 50600 36964
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 65656 36476 65720 36480
rect 65656 36420 65660 36476
rect 65660 36420 65716 36476
rect 65716 36420 65720 36476
rect 65656 36416 65720 36420
rect 65736 36476 65800 36480
rect 65736 36420 65740 36476
rect 65740 36420 65796 36476
rect 65796 36420 65800 36476
rect 65736 36416 65800 36420
rect 65816 36476 65880 36480
rect 65816 36420 65820 36476
rect 65820 36420 65876 36476
rect 65876 36420 65880 36476
rect 65816 36416 65880 36420
rect 65896 36476 65960 36480
rect 65896 36420 65900 36476
rect 65900 36420 65956 36476
rect 65956 36420 65960 36476
rect 65896 36416 65960 36420
rect 19576 35932 19640 35936
rect 19576 35876 19580 35932
rect 19580 35876 19636 35932
rect 19636 35876 19640 35932
rect 19576 35872 19640 35876
rect 19656 35932 19720 35936
rect 19656 35876 19660 35932
rect 19660 35876 19716 35932
rect 19716 35876 19720 35932
rect 19656 35872 19720 35876
rect 19736 35932 19800 35936
rect 19736 35876 19740 35932
rect 19740 35876 19796 35932
rect 19796 35876 19800 35932
rect 19736 35872 19800 35876
rect 19816 35932 19880 35936
rect 19816 35876 19820 35932
rect 19820 35876 19876 35932
rect 19876 35876 19880 35932
rect 19816 35872 19880 35876
rect 50296 35932 50360 35936
rect 50296 35876 50300 35932
rect 50300 35876 50356 35932
rect 50356 35876 50360 35932
rect 50296 35872 50360 35876
rect 50376 35932 50440 35936
rect 50376 35876 50380 35932
rect 50380 35876 50436 35932
rect 50436 35876 50440 35932
rect 50376 35872 50440 35876
rect 50456 35932 50520 35936
rect 50456 35876 50460 35932
rect 50460 35876 50516 35932
rect 50516 35876 50520 35932
rect 50456 35872 50520 35876
rect 50536 35932 50600 35936
rect 50536 35876 50540 35932
rect 50540 35876 50596 35932
rect 50596 35876 50600 35932
rect 50536 35872 50600 35876
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 65656 35388 65720 35392
rect 65656 35332 65660 35388
rect 65660 35332 65716 35388
rect 65716 35332 65720 35388
rect 65656 35328 65720 35332
rect 65736 35388 65800 35392
rect 65736 35332 65740 35388
rect 65740 35332 65796 35388
rect 65796 35332 65800 35388
rect 65736 35328 65800 35332
rect 65816 35388 65880 35392
rect 65816 35332 65820 35388
rect 65820 35332 65876 35388
rect 65876 35332 65880 35388
rect 65816 35328 65880 35332
rect 65896 35388 65960 35392
rect 65896 35332 65900 35388
rect 65900 35332 65956 35388
rect 65956 35332 65960 35388
rect 65896 35328 65960 35332
rect 19576 34844 19640 34848
rect 19576 34788 19580 34844
rect 19580 34788 19636 34844
rect 19636 34788 19640 34844
rect 19576 34784 19640 34788
rect 19656 34844 19720 34848
rect 19656 34788 19660 34844
rect 19660 34788 19716 34844
rect 19716 34788 19720 34844
rect 19656 34784 19720 34788
rect 19736 34844 19800 34848
rect 19736 34788 19740 34844
rect 19740 34788 19796 34844
rect 19796 34788 19800 34844
rect 19736 34784 19800 34788
rect 19816 34844 19880 34848
rect 19816 34788 19820 34844
rect 19820 34788 19876 34844
rect 19876 34788 19880 34844
rect 19816 34784 19880 34788
rect 50296 34844 50360 34848
rect 50296 34788 50300 34844
rect 50300 34788 50356 34844
rect 50356 34788 50360 34844
rect 50296 34784 50360 34788
rect 50376 34844 50440 34848
rect 50376 34788 50380 34844
rect 50380 34788 50436 34844
rect 50436 34788 50440 34844
rect 50376 34784 50440 34788
rect 50456 34844 50520 34848
rect 50456 34788 50460 34844
rect 50460 34788 50516 34844
rect 50516 34788 50520 34844
rect 50456 34784 50520 34788
rect 50536 34844 50600 34848
rect 50536 34788 50540 34844
rect 50540 34788 50596 34844
rect 50596 34788 50600 34844
rect 50536 34784 50600 34788
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 65656 34300 65720 34304
rect 65656 34244 65660 34300
rect 65660 34244 65716 34300
rect 65716 34244 65720 34300
rect 65656 34240 65720 34244
rect 65736 34300 65800 34304
rect 65736 34244 65740 34300
rect 65740 34244 65796 34300
rect 65796 34244 65800 34300
rect 65736 34240 65800 34244
rect 65816 34300 65880 34304
rect 65816 34244 65820 34300
rect 65820 34244 65876 34300
rect 65876 34244 65880 34300
rect 65816 34240 65880 34244
rect 65896 34300 65960 34304
rect 65896 34244 65900 34300
rect 65900 34244 65956 34300
rect 65956 34244 65960 34300
rect 65896 34240 65960 34244
rect 19576 33756 19640 33760
rect 19576 33700 19580 33756
rect 19580 33700 19636 33756
rect 19636 33700 19640 33756
rect 19576 33696 19640 33700
rect 19656 33756 19720 33760
rect 19656 33700 19660 33756
rect 19660 33700 19716 33756
rect 19716 33700 19720 33756
rect 19656 33696 19720 33700
rect 19736 33756 19800 33760
rect 19736 33700 19740 33756
rect 19740 33700 19796 33756
rect 19796 33700 19800 33756
rect 19736 33696 19800 33700
rect 19816 33756 19880 33760
rect 19816 33700 19820 33756
rect 19820 33700 19876 33756
rect 19876 33700 19880 33756
rect 19816 33696 19880 33700
rect 50296 33756 50360 33760
rect 50296 33700 50300 33756
rect 50300 33700 50356 33756
rect 50356 33700 50360 33756
rect 50296 33696 50360 33700
rect 50376 33756 50440 33760
rect 50376 33700 50380 33756
rect 50380 33700 50436 33756
rect 50436 33700 50440 33756
rect 50376 33696 50440 33700
rect 50456 33756 50520 33760
rect 50456 33700 50460 33756
rect 50460 33700 50516 33756
rect 50516 33700 50520 33756
rect 50456 33696 50520 33700
rect 50536 33756 50600 33760
rect 50536 33700 50540 33756
rect 50540 33700 50596 33756
rect 50596 33700 50600 33756
rect 50536 33696 50600 33700
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 65656 33212 65720 33216
rect 65656 33156 65660 33212
rect 65660 33156 65716 33212
rect 65716 33156 65720 33212
rect 65656 33152 65720 33156
rect 65736 33212 65800 33216
rect 65736 33156 65740 33212
rect 65740 33156 65796 33212
rect 65796 33156 65800 33212
rect 65736 33152 65800 33156
rect 65816 33212 65880 33216
rect 65816 33156 65820 33212
rect 65820 33156 65876 33212
rect 65876 33156 65880 33212
rect 65816 33152 65880 33156
rect 65896 33212 65960 33216
rect 65896 33156 65900 33212
rect 65900 33156 65956 33212
rect 65956 33156 65960 33212
rect 65896 33152 65960 33156
rect 19576 32668 19640 32672
rect 19576 32612 19580 32668
rect 19580 32612 19636 32668
rect 19636 32612 19640 32668
rect 19576 32608 19640 32612
rect 19656 32668 19720 32672
rect 19656 32612 19660 32668
rect 19660 32612 19716 32668
rect 19716 32612 19720 32668
rect 19656 32608 19720 32612
rect 19736 32668 19800 32672
rect 19736 32612 19740 32668
rect 19740 32612 19796 32668
rect 19796 32612 19800 32668
rect 19736 32608 19800 32612
rect 19816 32668 19880 32672
rect 19816 32612 19820 32668
rect 19820 32612 19876 32668
rect 19876 32612 19880 32668
rect 19816 32608 19880 32612
rect 50296 32668 50360 32672
rect 50296 32612 50300 32668
rect 50300 32612 50356 32668
rect 50356 32612 50360 32668
rect 50296 32608 50360 32612
rect 50376 32668 50440 32672
rect 50376 32612 50380 32668
rect 50380 32612 50436 32668
rect 50436 32612 50440 32668
rect 50376 32608 50440 32612
rect 50456 32668 50520 32672
rect 50456 32612 50460 32668
rect 50460 32612 50516 32668
rect 50516 32612 50520 32668
rect 50456 32608 50520 32612
rect 50536 32668 50600 32672
rect 50536 32612 50540 32668
rect 50540 32612 50596 32668
rect 50596 32612 50600 32668
rect 50536 32608 50600 32612
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 65656 32124 65720 32128
rect 65656 32068 65660 32124
rect 65660 32068 65716 32124
rect 65716 32068 65720 32124
rect 65656 32064 65720 32068
rect 65736 32124 65800 32128
rect 65736 32068 65740 32124
rect 65740 32068 65796 32124
rect 65796 32068 65800 32124
rect 65736 32064 65800 32068
rect 65816 32124 65880 32128
rect 65816 32068 65820 32124
rect 65820 32068 65876 32124
rect 65876 32068 65880 32124
rect 65816 32064 65880 32068
rect 65896 32124 65960 32128
rect 65896 32068 65900 32124
rect 65900 32068 65956 32124
rect 65956 32068 65960 32124
rect 65896 32064 65960 32068
rect 19576 31580 19640 31584
rect 19576 31524 19580 31580
rect 19580 31524 19636 31580
rect 19636 31524 19640 31580
rect 19576 31520 19640 31524
rect 19656 31580 19720 31584
rect 19656 31524 19660 31580
rect 19660 31524 19716 31580
rect 19716 31524 19720 31580
rect 19656 31520 19720 31524
rect 19736 31580 19800 31584
rect 19736 31524 19740 31580
rect 19740 31524 19796 31580
rect 19796 31524 19800 31580
rect 19736 31520 19800 31524
rect 19816 31580 19880 31584
rect 19816 31524 19820 31580
rect 19820 31524 19876 31580
rect 19876 31524 19880 31580
rect 19816 31520 19880 31524
rect 50296 31580 50360 31584
rect 50296 31524 50300 31580
rect 50300 31524 50356 31580
rect 50356 31524 50360 31580
rect 50296 31520 50360 31524
rect 50376 31580 50440 31584
rect 50376 31524 50380 31580
rect 50380 31524 50436 31580
rect 50436 31524 50440 31580
rect 50376 31520 50440 31524
rect 50456 31580 50520 31584
rect 50456 31524 50460 31580
rect 50460 31524 50516 31580
rect 50516 31524 50520 31580
rect 50456 31520 50520 31524
rect 50536 31580 50600 31584
rect 50536 31524 50540 31580
rect 50540 31524 50596 31580
rect 50596 31524 50600 31580
rect 50536 31520 50600 31524
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 65656 31036 65720 31040
rect 65656 30980 65660 31036
rect 65660 30980 65716 31036
rect 65716 30980 65720 31036
rect 65656 30976 65720 30980
rect 65736 31036 65800 31040
rect 65736 30980 65740 31036
rect 65740 30980 65796 31036
rect 65796 30980 65800 31036
rect 65736 30976 65800 30980
rect 65816 31036 65880 31040
rect 65816 30980 65820 31036
rect 65820 30980 65876 31036
rect 65876 30980 65880 31036
rect 65816 30976 65880 30980
rect 65896 31036 65960 31040
rect 65896 30980 65900 31036
rect 65900 30980 65956 31036
rect 65956 30980 65960 31036
rect 65896 30976 65960 30980
rect 19576 30492 19640 30496
rect 19576 30436 19580 30492
rect 19580 30436 19636 30492
rect 19636 30436 19640 30492
rect 19576 30432 19640 30436
rect 19656 30492 19720 30496
rect 19656 30436 19660 30492
rect 19660 30436 19716 30492
rect 19716 30436 19720 30492
rect 19656 30432 19720 30436
rect 19736 30492 19800 30496
rect 19736 30436 19740 30492
rect 19740 30436 19796 30492
rect 19796 30436 19800 30492
rect 19736 30432 19800 30436
rect 19816 30492 19880 30496
rect 19816 30436 19820 30492
rect 19820 30436 19876 30492
rect 19876 30436 19880 30492
rect 19816 30432 19880 30436
rect 50296 30492 50360 30496
rect 50296 30436 50300 30492
rect 50300 30436 50356 30492
rect 50356 30436 50360 30492
rect 50296 30432 50360 30436
rect 50376 30492 50440 30496
rect 50376 30436 50380 30492
rect 50380 30436 50436 30492
rect 50436 30436 50440 30492
rect 50376 30432 50440 30436
rect 50456 30492 50520 30496
rect 50456 30436 50460 30492
rect 50460 30436 50516 30492
rect 50516 30436 50520 30492
rect 50456 30432 50520 30436
rect 50536 30492 50600 30496
rect 50536 30436 50540 30492
rect 50540 30436 50596 30492
rect 50596 30436 50600 30492
rect 50536 30432 50600 30436
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 65656 29948 65720 29952
rect 65656 29892 65660 29948
rect 65660 29892 65716 29948
rect 65716 29892 65720 29948
rect 65656 29888 65720 29892
rect 65736 29948 65800 29952
rect 65736 29892 65740 29948
rect 65740 29892 65796 29948
rect 65796 29892 65800 29948
rect 65736 29888 65800 29892
rect 65816 29948 65880 29952
rect 65816 29892 65820 29948
rect 65820 29892 65876 29948
rect 65876 29892 65880 29948
rect 65816 29888 65880 29892
rect 65896 29948 65960 29952
rect 65896 29892 65900 29948
rect 65900 29892 65956 29948
rect 65956 29892 65960 29948
rect 65896 29888 65960 29892
rect 19576 29404 19640 29408
rect 19576 29348 19580 29404
rect 19580 29348 19636 29404
rect 19636 29348 19640 29404
rect 19576 29344 19640 29348
rect 19656 29404 19720 29408
rect 19656 29348 19660 29404
rect 19660 29348 19716 29404
rect 19716 29348 19720 29404
rect 19656 29344 19720 29348
rect 19736 29404 19800 29408
rect 19736 29348 19740 29404
rect 19740 29348 19796 29404
rect 19796 29348 19800 29404
rect 19736 29344 19800 29348
rect 19816 29404 19880 29408
rect 19816 29348 19820 29404
rect 19820 29348 19876 29404
rect 19876 29348 19880 29404
rect 19816 29344 19880 29348
rect 50296 29404 50360 29408
rect 50296 29348 50300 29404
rect 50300 29348 50356 29404
rect 50356 29348 50360 29404
rect 50296 29344 50360 29348
rect 50376 29404 50440 29408
rect 50376 29348 50380 29404
rect 50380 29348 50436 29404
rect 50436 29348 50440 29404
rect 50376 29344 50440 29348
rect 50456 29404 50520 29408
rect 50456 29348 50460 29404
rect 50460 29348 50516 29404
rect 50516 29348 50520 29404
rect 50456 29344 50520 29348
rect 50536 29404 50600 29408
rect 50536 29348 50540 29404
rect 50540 29348 50596 29404
rect 50596 29348 50600 29404
rect 50536 29344 50600 29348
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 65656 28860 65720 28864
rect 65656 28804 65660 28860
rect 65660 28804 65716 28860
rect 65716 28804 65720 28860
rect 65656 28800 65720 28804
rect 65736 28860 65800 28864
rect 65736 28804 65740 28860
rect 65740 28804 65796 28860
rect 65796 28804 65800 28860
rect 65736 28800 65800 28804
rect 65816 28860 65880 28864
rect 65816 28804 65820 28860
rect 65820 28804 65876 28860
rect 65876 28804 65880 28860
rect 65816 28800 65880 28804
rect 65896 28860 65960 28864
rect 65896 28804 65900 28860
rect 65900 28804 65956 28860
rect 65956 28804 65960 28860
rect 65896 28800 65960 28804
rect 19576 28316 19640 28320
rect 19576 28260 19580 28316
rect 19580 28260 19636 28316
rect 19636 28260 19640 28316
rect 19576 28256 19640 28260
rect 19656 28316 19720 28320
rect 19656 28260 19660 28316
rect 19660 28260 19716 28316
rect 19716 28260 19720 28316
rect 19656 28256 19720 28260
rect 19736 28316 19800 28320
rect 19736 28260 19740 28316
rect 19740 28260 19796 28316
rect 19796 28260 19800 28316
rect 19736 28256 19800 28260
rect 19816 28316 19880 28320
rect 19816 28260 19820 28316
rect 19820 28260 19876 28316
rect 19876 28260 19880 28316
rect 19816 28256 19880 28260
rect 50296 28316 50360 28320
rect 50296 28260 50300 28316
rect 50300 28260 50356 28316
rect 50356 28260 50360 28316
rect 50296 28256 50360 28260
rect 50376 28316 50440 28320
rect 50376 28260 50380 28316
rect 50380 28260 50436 28316
rect 50436 28260 50440 28316
rect 50376 28256 50440 28260
rect 50456 28316 50520 28320
rect 50456 28260 50460 28316
rect 50460 28260 50516 28316
rect 50516 28260 50520 28316
rect 50456 28256 50520 28260
rect 50536 28316 50600 28320
rect 50536 28260 50540 28316
rect 50540 28260 50596 28316
rect 50596 28260 50600 28316
rect 50536 28256 50600 28260
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 65656 27772 65720 27776
rect 65656 27716 65660 27772
rect 65660 27716 65716 27772
rect 65716 27716 65720 27772
rect 65656 27712 65720 27716
rect 65736 27772 65800 27776
rect 65736 27716 65740 27772
rect 65740 27716 65796 27772
rect 65796 27716 65800 27772
rect 65736 27712 65800 27716
rect 65816 27772 65880 27776
rect 65816 27716 65820 27772
rect 65820 27716 65876 27772
rect 65876 27716 65880 27772
rect 65816 27712 65880 27716
rect 65896 27772 65960 27776
rect 65896 27716 65900 27772
rect 65900 27716 65956 27772
rect 65956 27716 65960 27772
rect 65896 27712 65960 27716
rect 19576 27228 19640 27232
rect 19576 27172 19580 27228
rect 19580 27172 19636 27228
rect 19636 27172 19640 27228
rect 19576 27168 19640 27172
rect 19656 27228 19720 27232
rect 19656 27172 19660 27228
rect 19660 27172 19716 27228
rect 19716 27172 19720 27228
rect 19656 27168 19720 27172
rect 19736 27228 19800 27232
rect 19736 27172 19740 27228
rect 19740 27172 19796 27228
rect 19796 27172 19800 27228
rect 19736 27168 19800 27172
rect 19816 27228 19880 27232
rect 19816 27172 19820 27228
rect 19820 27172 19876 27228
rect 19876 27172 19880 27228
rect 19816 27168 19880 27172
rect 50296 27228 50360 27232
rect 50296 27172 50300 27228
rect 50300 27172 50356 27228
rect 50356 27172 50360 27228
rect 50296 27168 50360 27172
rect 50376 27228 50440 27232
rect 50376 27172 50380 27228
rect 50380 27172 50436 27228
rect 50436 27172 50440 27228
rect 50376 27168 50440 27172
rect 50456 27228 50520 27232
rect 50456 27172 50460 27228
rect 50460 27172 50516 27228
rect 50516 27172 50520 27228
rect 50456 27168 50520 27172
rect 50536 27228 50600 27232
rect 50536 27172 50540 27228
rect 50540 27172 50596 27228
rect 50596 27172 50600 27228
rect 50536 27168 50600 27172
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 65656 26684 65720 26688
rect 65656 26628 65660 26684
rect 65660 26628 65716 26684
rect 65716 26628 65720 26684
rect 65656 26624 65720 26628
rect 65736 26684 65800 26688
rect 65736 26628 65740 26684
rect 65740 26628 65796 26684
rect 65796 26628 65800 26684
rect 65736 26624 65800 26628
rect 65816 26684 65880 26688
rect 65816 26628 65820 26684
rect 65820 26628 65876 26684
rect 65876 26628 65880 26684
rect 65816 26624 65880 26628
rect 65896 26684 65960 26688
rect 65896 26628 65900 26684
rect 65900 26628 65956 26684
rect 65956 26628 65960 26684
rect 65896 26624 65960 26628
rect 19576 26140 19640 26144
rect 19576 26084 19580 26140
rect 19580 26084 19636 26140
rect 19636 26084 19640 26140
rect 19576 26080 19640 26084
rect 19656 26140 19720 26144
rect 19656 26084 19660 26140
rect 19660 26084 19716 26140
rect 19716 26084 19720 26140
rect 19656 26080 19720 26084
rect 19736 26140 19800 26144
rect 19736 26084 19740 26140
rect 19740 26084 19796 26140
rect 19796 26084 19800 26140
rect 19736 26080 19800 26084
rect 19816 26140 19880 26144
rect 19816 26084 19820 26140
rect 19820 26084 19876 26140
rect 19876 26084 19880 26140
rect 19816 26080 19880 26084
rect 50296 26140 50360 26144
rect 50296 26084 50300 26140
rect 50300 26084 50356 26140
rect 50356 26084 50360 26140
rect 50296 26080 50360 26084
rect 50376 26140 50440 26144
rect 50376 26084 50380 26140
rect 50380 26084 50436 26140
rect 50436 26084 50440 26140
rect 50376 26080 50440 26084
rect 50456 26140 50520 26144
rect 50456 26084 50460 26140
rect 50460 26084 50516 26140
rect 50516 26084 50520 26140
rect 50456 26080 50520 26084
rect 50536 26140 50600 26144
rect 50536 26084 50540 26140
rect 50540 26084 50596 26140
rect 50596 26084 50600 26140
rect 50536 26080 50600 26084
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 65656 25596 65720 25600
rect 65656 25540 65660 25596
rect 65660 25540 65716 25596
rect 65716 25540 65720 25596
rect 65656 25536 65720 25540
rect 65736 25596 65800 25600
rect 65736 25540 65740 25596
rect 65740 25540 65796 25596
rect 65796 25540 65800 25596
rect 65736 25536 65800 25540
rect 65816 25596 65880 25600
rect 65816 25540 65820 25596
rect 65820 25540 65876 25596
rect 65876 25540 65880 25596
rect 65816 25536 65880 25540
rect 65896 25596 65960 25600
rect 65896 25540 65900 25596
rect 65900 25540 65956 25596
rect 65956 25540 65960 25596
rect 65896 25536 65960 25540
rect 19576 25052 19640 25056
rect 19576 24996 19580 25052
rect 19580 24996 19636 25052
rect 19636 24996 19640 25052
rect 19576 24992 19640 24996
rect 19656 25052 19720 25056
rect 19656 24996 19660 25052
rect 19660 24996 19716 25052
rect 19716 24996 19720 25052
rect 19656 24992 19720 24996
rect 19736 25052 19800 25056
rect 19736 24996 19740 25052
rect 19740 24996 19796 25052
rect 19796 24996 19800 25052
rect 19736 24992 19800 24996
rect 19816 25052 19880 25056
rect 19816 24996 19820 25052
rect 19820 24996 19876 25052
rect 19876 24996 19880 25052
rect 19816 24992 19880 24996
rect 50296 25052 50360 25056
rect 50296 24996 50300 25052
rect 50300 24996 50356 25052
rect 50356 24996 50360 25052
rect 50296 24992 50360 24996
rect 50376 25052 50440 25056
rect 50376 24996 50380 25052
rect 50380 24996 50436 25052
rect 50436 24996 50440 25052
rect 50376 24992 50440 24996
rect 50456 25052 50520 25056
rect 50456 24996 50460 25052
rect 50460 24996 50516 25052
rect 50516 24996 50520 25052
rect 50456 24992 50520 24996
rect 50536 25052 50600 25056
rect 50536 24996 50540 25052
rect 50540 24996 50596 25052
rect 50596 24996 50600 25052
rect 50536 24992 50600 24996
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 65656 24508 65720 24512
rect 65656 24452 65660 24508
rect 65660 24452 65716 24508
rect 65716 24452 65720 24508
rect 65656 24448 65720 24452
rect 65736 24508 65800 24512
rect 65736 24452 65740 24508
rect 65740 24452 65796 24508
rect 65796 24452 65800 24508
rect 65736 24448 65800 24452
rect 65816 24508 65880 24512
rect 65816 24452 65820 24508
rect 65820 24452 65876 24508
rect 65876 24452 65880 24508
rect 65816 24448 65880 24452
rect 65896 24508 65960 24512
rect 65896 24452 65900 24508
rect 65900 24452 65956 24508
rect 65956 24452 65960 24508
rect 65896 24448 65960 24452
rect 19576 23964 19640 23968
rect 19576 23908 19580 23964
rect 19580 23908 19636 23964
rect 19636 23908 19640 23964
rect 19576 23904 19640 23908
rect 19656 23964 19720 23968
rect 19656 23908 19660 23964
rect 19660 23908 19716 23964
rect 19716 23908 19720 23964
rect 19656 23904 19720 23908
rect 19736 23964 19800 23968
rect 19736 23908 19740 23964
rect 19740 23908 19796 23964
rect 19796 23908 19800 23964
rect 19736 23904 19800 23908
rect 19816 23964 19880 23968
rect 19816 23908 19820 23964
rect 19820 23908 19876 23964
rect 19876 23908 19880 23964
rect 19816 23904 19880 23908
rect 50296 23964 50360 23968
rect 50296 23908 50300 23964
rect 50300 23908 50356 23964
rect 50356 23908 50360 23964
rect 50296 23904 50360 23908
rect 50376 23964 50440 23968
rect 50376 23908 50380 23964
rect 50380 23908 50436 23964
rect 50436 23908 50440 23964
rect 50376 23904 50440 23908
rect 50456 23964 50520 23968
rect 50456 23908 50460 23964
rect 50460 23908 50516 23964
rect 50516 23908 50520 23964
rect 50456 23904 50520 23908
rect 50536 23964 50600 23968
rect 50536 23908 50540 23964
rect 50540 23908 50596 23964
rect 50596 23908 50600 23964
rect 50536 23904 50600 23908
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 65656 23420 65720 23424
rect 65656 23364 65660 23420
rect 65660 23364 65716 23420
rect 65716 23364 65720 23420
rect 65656 23360 65720 23364
rect 65736 23420 65800 23424
rect 65736 23364 65740 23420
rect 65740 23364 65796 23420
rect 65796 23364 65800 23420
rect 65736 23360 65800 23364
rect 65816 23420 65880 23424
rect 65816 23364 65820 23420
rect 65820 23364 65876 23420
rect 65876 23364 65880 23420
rect 65816 23360 65880 23364
rect 65896 23420 65960 23424
rect 65896 23364 65900 23420
rect 65900 23364 65956 23420
rect 65956 23364 65960 23420
rect 65896 23360 65960 23364
rect 19576 22876 19640 22880
rect 19576 22820 19580 22876
rect 19580 22820 19636 22876
rect 19636 22820 19640 22876
rect 19576 22816 19640 22820
rect 19656 22876 19720 22880
rect 19656 22820 19660 22876
rect 19660 22820 19716 22876
rect 19716 22820 19720 22876
rect 19656 22816 19720 22820
rect 19736 22876 19800 22880
rect 19736 22820 19740 22876
rect 19740 22820 19796 22876
rect 19796 22820 19800 22876
rect 19736 22816 19800 22820
rect 19816 22876 19880 22880
rect 19816 22820 19820 22876
rect 19820 22820 19876 22876
rect 19876 22820 19880 22876
rect 19816 22816 19880 22820
rect 50296 22876 50360 22880
rect 50296 22820 50300 22876
rect 50300 22820 50356 22876
rect 50356 22820 50360 22876
rect 50296 22816 50360 22820
rect 50376 22876 50440 22880
rect 50376 22820 50380 22876
rect 50380 22820 50436 22876
rect 50436 22820 50440 22876
rect 50376 22816 50440 22820
rect 50456 22876 50520 22880
rect 50456 22820 50460 22876
rect 50460 22820 50516 22876
rect 50516 22820 50520 22876
rect 50456 22816 50520 22820
rect 50536 22876 50600 22880
rect 50536 22820 50540 22876
rect 50540 22820 50596 22876
rect 50596 22820 50600 22876
rect 50536 22816 50600 22820
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 65656 22332 65720 22336
rect 65656 22276 65660 22332
rect 65660 22276 65716 22332
rect 65716 22276 65720 22332
rect 65656 22272 65720 22276
rect 65736 22332 65800 22336
rect 65736 22276 65740 22332
rect 65740 22276 65796 22332
rect 65796 22276 65800 22332
rect 65736 22272 65800 22276
rect 65816 22332 65880 22336
rect 65816 22276 65820 22332
rect 65820 22276 65876 22332
rect 65876 22276 65880 22332
rect 65816 22272 65880 22276
rect 65896 22332 65960 22336
rect 65896 22276 65900 22332
rect 65900 22276 65956 22332
rect 65956 22276 65960 22332
rect 65896 22272 65960 22276
rect 19576 21788 19640 21792
rect 19576 21732 19580 21788
rect 19580 21732 19636 21788
rect 19636 21732 19640 21788
rect 19576 21728 19640 21732
rect 19656 21788 19720 21792
rect 19656 21732 19660 21788
rect 19660 21732 19716 21788
rect 19716 21732 19720 21788
rect 19656 21728 19720 21732
rect 19736 21788 19800 21792
rect 19736 21732 19740 21788
rect 19740 21732 19796 21788
rect 19796 21732 19800 21788
rect 19736 21728 19800 21732
rect 19816 21788 19880 21792
rect 19816 21732 19820 21788
rect 19820 21732 19876 21788
rect 19876 21732 19880 21788
rect 19816 21728 19880 21732
rect 50296 21788 50360 21792
rect 50296 21732 50300 21788
rect 50300 21732 50356 21788
rect 50356 21732 50360 21788
rect 50296 21728 50360 21732
rect 50376 21788 50440 21792
rect 50376 21732 50380 21788
rect 50380 21732 50436 21788
rect 50436 21732 50440 21788
rect 50376 21728 50440 21732
rect 50456 21788 50520 21792
rect 50456 21732 50460 21788
rect 50460 21732 50516 21788
rect 50516 21732 50520 21788
rect 50456 21728 50520 21732
rect 50536 21788 50600 21792
rect 50536 21732 50540 21788
rect 50540 21732 50596 21788
rect 50596 21732 50600 21788
rect 50536 21728 50600 21732
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 65656 21244 65720 21248
rect 65656 21188 65660 21244
rect 65660 21188 65716 21244
rect 65716 21188 65720 21244
rect 65656 21184 65720 21188
rect 65736 21244 65800 21248
rect 65736 21188 65740 21244
rect 65740 21188 65796 21244
rect 65796 21188 65800 21244
rect 65736 21184 65800 21188
rect 65816 21244 65880 21248
rect 65816 21188 65820 21244
rect 65820 21188 65876 21244
rect 65876 21188 65880 21244
rect 65816 21184 65880 21188
rect 65896 21244 65960 21248
rect 65896 21188 65900 21244
rect 65900 21188 65956 21244
rect 65956 21188 65960 21244
rect 65896 21184 65960 21188
rect 19576 20700 19640 20704
rect 19576 20644 19580 20700
rect 19580 20644 19636 20700
rect 19636 20644 19640 20700
rect 19576 20640 19640 20644
rect 19656 20700 19720 20704
rect 19656 20644 19660 20700
rect 19660 20644 19716 20700
rect 19716 20644 19720 20700
rect 19656 20640 19720 20644
rect 19736 20700 19800 20704
rect 19736 20644 19740 20700
rect 19740 20644 19796 20700
rect 19796 20644 19800 20700
rect 19736 20640 19800 20644
rect 19816 20700 19880 20704
rect 19816 20644 19820 20700
rect 19820 20644 19876 20700
rect 19876 20644 19880 20700
rect 19816 20640 19880 20644
rect 50296 20700 50360 20704
rect 50296 20644 50300 20700
rect 50300 20644 50356 20700
rect 50356 20644 50360 20700
rect 50296 20640 50360 20644
rect 50376 20700 50440 20704
rect 50376 20644 50380 20700
rect 50380 20644 50436 20700
rect 50436 20644 50440 20700
rect 50376 20640 50440 20644
rect 50456 20700 50520 20704
rect 50456 20644 50460 20700
rect 50460 20644 50516 20700
rect 50516 20644 50520 20700
rect 50456 20640 50520 20644
rect 50536 20700 50600 20704
rect 50536 20644 50540 20700
rect 50540 20644 50596 20700
rect 50596 20644 50600 20700
rect 50536 20640 50600 20644
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 65656 20156 65720 20160
rect 65656 20100 65660 20156
rect 65660 20100 65716 20156
rect 65716 20100 65720 20156
rect 65656 20096 65720 20100
rect 65736 20156 65800 20160
rect 65736 20100 65740 20156
rect 65740 20100 65796 20156
rect 65796 20100 65800 20156
rect 65736 20096 65800 20100
rect 65816 20156 65880 20160
rect 65816 20100 65820 20156
rect 65820 20100 65876 20156
rect 65876 20100 65880 20156
rect 65816 20096 65880 20100
rect 65896 20156 65960 20160
rect 65896 20100 65900 20156
rect 65900 20100 65956 20156
rect 65956 20100 65960 20156
rect 65896 20096 65960 20100
rect 19576 19612 19640 19616
rect 19576 19556 19580 19612
rect 19580 19556 19636 19612
rect 19636 19556 19640 19612
rect 19576 19552 19640 19556
rect 19656 19612 19720 19616
rect 19656 19556 19660 19612
rect 19660 19556 19716 19612
rect 19716 19556 19720 19612
rect 19656 19552 19720 19556
rect 19736 19612 19800 19616
rect 19736 19556 19740 19612
rect 19740 19556 19796 19612
rect 19796 19556 19800 19612
rect 19736 19552 19800 19556
rect 19816 19612 19880 19616
rect 19816 19556 19820 19612
rect 19820 19556 19876 19612
rect 19876 19556 19880 19612
rect 19816 19552 19880 19556
rect 50296 19612 50360 19616
rect 50296 19556 50300 19612
rect 50300 19556 50356 19612
rect 50356 19556 50360 19612
rect 50296 19552 50360 19556
rect 50376 19612 50440 19616
rect 50376 19556 50380 19612
rect 50380 19556 50436 19612
rect 50436 19556 50440 19612
rect 50376 19552 50440 19556
rect 50456 19612 50520 19616
rect 50456 19556 50460 19612
rect 50460 19556 50516 19612
rect 50516 19556 50520 19612
rect 50456 19552 50520 19556
rect 50536 19612 50600 19616
rect 50536 19556 50540 19612
rect 50540 19556 50596 19612
rect 50596 19556 50600 19612
rect 50536 19552 50600 19556
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 65656 19068 65720 19072
rect 65656 19012 65660 19068
rect 65660 19012 65716 19068
rect 65716 19012 65720 19068
rect 65656 19008 65720 19012
rect 65736 19068 65800 19072
rect 65736 19012 65740 19068
rect 65740 19012 65796 19068
rect 65796 19012 65800 19068
rect 65736 19008 65800 19012
rect 65816 19068 65880 19072
rect 65816 19012 65820 19068
rect 65820 19012 65876 19068
rect 65876 19012 65880 19068
rect 65816 19008 65880 19012
rect 65896 19068 65960 19072
rect 65896 19012 65900 19068
rect 65900 19012 65956 19068
rect 65956 19012 65960 19068
rect 65896 19008 65960 19012
rect 19576 18524 19640 18528
rect 19576 18468 19580 18524
rect 19580 18468 19636 18524
rect 19636 18468 19640 18524
rect 19576 18464 19640 18468
rect 19656 18524 19720 18528
rect 19656 18468 19660 18524
rect 19660 18468 19716 18524
rect 19716 18468 19720 18524
rect 19656 18464 19720 18468
rect 19736 18524 19800 18528
rect 19736 18468 19740 18524
rect 19740 18468 19796 18524
rect 19796 18468 19800 18524
rect 19736 18464 19800 18468
rect 19816 18524 19880 18528
rect 19816 18468 19820 18524
rect 19820 18468 19876 18524
rect 19876 18468 19880 18524
rect 19816 18464 19880 18468
rect 50296 18524 50360 18528
rect 50296 18468 50300 18524
rect 50300 18468 50356 18524
rect 50356 18468 50360 18524
rect 50296 18464 50360 18468
rect 50376 18524 50440 18528
rect 50376 18468 50380 18524
rect 50380 18468 50436 18524
rect 50436 18468 50440 18524
rect 50376 18464 50440 18468
rect 50456 18524 50520 18528
rect 50456 18468 50460 18524
rect 50460 18468 50516 18524
rect 50516 18468 50520 18524
rect 50456 18464 50520 18468
rect 50536 18524 50600 18528
rect 50536 18468 50540 18524
rect 50540 18468 50596 18524
rect 50596 18468 50600 18524
rect 50536 18464 50600 18468
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 65656 17980 65720 17984
rect 65656 17924 65660 17980
rect 65660 17924 65716 17980
rect 65716 17924 65720 17980
rect 65656 17920 65720 17924
rect 65736 17980 65800 17984
rect 65736 17924 65740 17980
rect 65740 17924 65796 17980
rect 65796 17924 65800 17980
rect 65736 17920 65800 17924
rect 65816 17980 65880 17984
rect 65816 17924 65820 17980
rect 65820 17924 65876 17980
rect 65876 17924 65880 17980
rect 65816 17920 65880 17924
rect 65896 17980 65960 17984
rect 65896 17924 65900 17980
rect 65900 17924 65956 17980
rect 65956 17924 65960 17980
rect 65896 17920 65960 17924
rect 19576 17436 19640 17440
rect 19576 17380 19580 17436
rect 19580 17380 19636 17436
rect 19636 17380 19640 17436
rect 19576 17376 19640 17380
rect 19656 17436 19720 17440
rect 19656 17380 19660 17436
rect 19660 17380 19716 17436
rect 19716 17380 19720 17436
rect 19656 17376 19720 17380
rect 19736 17436 19800 17440
rect 19736 17380 19740 17436
rect 19740 17380 19796 17436
rect 19796 17380 19800 17436
rect 19736 17376 19800 17380
rect 19816 17436 19880 17440
rect 19816 17380 19820 17436
rect 19820 17380 19876 17436
rect 19876 17380 19880 17436
rect 19816 17376 19880 17380
rect 50296 17436 50360 17440
rect 50296 17380 50300 17436
rect 50300 17380 50356 17436
rect 50356 17380 50360 17436
rect 50296 17376 50360 17380
rect 50376 17436 50440 17440
rect 50376 17380 50380 17436
rect 50380 17380 50436 17436
rect 50436 17380 50440 17436
rect 50376 17376 50440 17380
rect 50456 17436 50520 17440
rect 50456 17380 50460 17436
rect 50460 17380 50516 17436
rect 50516 17380 50520 17436
rect 50456 17376 50520 17380
rect 50536 17436 50600 17440
rect 50536 17380 50540 17436
rect 50540 17380 50596 17436
rect 50596 17380 50600 17436
rect 50536 17376 50600 17380
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 65656 16892 65720 16896
rect 65656 16836 65660 16892
rect 65660 16836 65716 16892
rect 65716 16836 65720 16892
rect 65656 16832 65720 16836
rect 65736 16892 65800 16896
rect 65736 16836 65740 16892
rect 65740 16836 65796 16892
rect 65796 16836 65800 16892
rect 65736 16832 65800 16836
rect 65816 16892 65880 16896
rect 65816 16836 65820 16892
rect 65820 16836 65876 16892
rect 65876 16836 65880 16892
rect 65816 16832 65880 16836
rect 65896 16892 65960 16896
rect 65896 16836 65900 16892
rect 65900 16836 65956 16892
rect 65956 16836 65960 16892
rect 65896 16832 65960 16836
rect 19576 16348 19640 16352
rect 19576 16292 19580 16348
rect 19580 16292 19636 16348
rect 19636 16292 19640 16348
rect 19576 16288 19640 16292
rect 19656 16348 19720 16352
rect 19656 16292 19660 16348
rect 19660 16292 19716 16348
rect 19716 16292 19720 16348
rect 19656 16288 19720 16292
rect 19736 16348 19800 16352
rect 19736 16292 19740 16348
rect 19740 16292 19796 16348
rect 19796 16292 19800 16348
rect 19736 16288 19800 16292
rect 19816 16348 19880 16352
rect 19816 16292 19820 16348
rect 19820 16292 19876 16348
rect 19876 16292 19880 16348
rect 19816 16288 19880 16292
rect 50296 16348 50360 16352
rect 50296 16292 50300 16348
rect 50300 16292 50356 16348
rect 50356 16292 50360 16348
rect 50296 16288 50360 16292
rect 50376 16348 50440 16352
rect 50376 16292 50380 16348
rect 50380 16292 50436 16348
rect 50436 16292 50440 16348
rect 50376 16288 50440 16292
rect 50456 16348 50520 16352
rect 50456 16292 50460 16348
rect 50460 16292 50516 16348
rect 50516 16292 50520 16348
rect 50456 16288 50520 16292
rect 50536 16348 50600 16352
rect 50536 16292 50540 16348
rect 50540 16292 50596 16348
rect 50596 16292 50600 16348
rect 50536 16288 50600 16292
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 65656 15804 65720 15808
rect 65656 15748 65660 15804
rect 65660 15748 65716 15804
rect 65716 15748 65720 15804
rect 65656 15744 65720 15748
rect 65736 15804 65800 15808
rect 65736 15748 65740 15804
rect 65740 15748 65796 15804
rect 65796 15748 65800 15804
rect 65736 15744 65800 15748
rect 65816 15804 65880 15808
rect 65816 15748 65820 15804
rect 65820 15748 65876 15804
rect 65876 15748 65880 15804
rect 65816 15744 65880 15748
rect 65896 15804 65960 15808
rect 65896 15748 65900 15804
rect 65900 15748 65956 15804
rect 65956 15748 65960 15804
rect 65896 15744 65960 15748
rect 19576 15260 19640 15264
rect 19576 15204 19580 15260
rect 19580 15204 19636 15260
rect 19636 15204 19640 15260
rect 19576 15200 19640 15204
rect 19656 15260 19720 15264
rect 19656 15204 19660 15260
rect 19660 15204 19716 15260
rect 19716 15204 19720 15260
rect 19656 15200 19720 15204
rect 19736 15260 19800 15264
rect 19736 15204 19740 15260
rect 19740 15204 19796 15260
rect 19796 15204 19800 15260
rect 19736 15200 19800 15204
rect 19816 15260 19880 15264
rect 19816 15204 19820 15260
rect 19820 15204 19876 15260
rect 19876 15204 19880 15260
rect 19816 15200 19880 15204
rect 50296 15260 50360 15264
rect 50296 15204 50300 15260
rect 50300 15204 50356 15260
rect 50356 15204 50360 15260
rect 50296 15200 50360 15204
rect 50376 15260 50440 15264
rect 50376 15204 50380 15260
rect 50380 15204 50436 15260
rect 50436 15204 50440 15260
rect 50376 15200 50440 15204
rect 50456 15260 50520 15264
rect 50456 15204 50460 15260
rect 50460 15204 50516 15260
rect 50516 15204 50520 15260
rect 50456 15200 50520 15204
rect 50536 15260 50600 15264
rect 50536 15204 50540 15260
rect 50540 15204 50596 15260
rect 50596 15204 50600 15260
rect 50536 15200 50600 15204
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 65656 14716 65720 14720
rect 65656 14660 65660 14716
rect 65660 14660 65716 14716
rect 65716 14660 65720 14716
rect 65656 14656 65720 14660
rect 65736 14716 65800 14720
rect 65736 14660 65740 14716
rect 65740 14660 65796 14716
rect 65796 14660 65800 14716
rect 65736 14656 65800 14660
rect 65816 14716 65880 14720
rect 65816 14660 65820 14716
rect 65820 14660 65876 14716
rect 65876 14660 65880 14716
rect 65816 14656 65880 14660
rect 65896 14716 65960 14720
rect 65896 14660 65900 14716
rect 65900 14660 65956 14716
rect 65956 14660 65960 14716
rect 65896 14656 65960 14660
rect 19576 14172 19640 14176
rect 19576 14116 19580 14172
rect 19580 14116 19636 14172
rect 19636 14116 19640 14172
rect 19576 14112 19640 14116
rect 19656 14172 19720 14176
rect 19656 14116 19660 14172
rect 19660 14116 19716 14172
rect 19716 14116 19720 14172
rect 19656 14112 19720 14116
rect 19736 14172 19800 14176
rect 19736 14116 19740 14172
rect 19740 14116 19796 14172
rect 19796 14116 19800 14172
rect 19736 14112 19800 14116
rect 19816 14172 19880 14176
rect 19816 14116 19820 14172
rect 19820 14116 19876 14172
rect 19876 14116 19880 14172
rect 19816 14112 19880 14116
rect 50296 14172 50360 14176
rect 50296 14116 50300 14172
rect 50300 14116 50356 14172
rect 50356 14116 50360 14172
rect 50296 14112 50360 14116
rect 50376 14172 50440 14176
rect 50376 14116 50380 14172
rect 50380 14116 50436 14172
rect 50436 14116 50440 14172
rect 50376 14112 50440 14116
rect 50456 14172 50520 14176
rect 50456 14116 50460 14172
rect 50460 14116 50516 14172
rect 50516 14116 50520 14172
rect 50456 14112 50520 14116
rect 50536 14172 50600 14176
rect 50536 14116 50540 14172
rect 50540 14116 50596 14172
rect 50596 14116 50600 14172
rect 50536 14112 50600 14116
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 65656 13628 65720 13632
rect 65656 13572 65660 13628
rect 65660 13572 65716 13628
rect 65716 13572 65720 13628
rect 65656 13568 65720 13572
rect 65736 13628 65800 13632
rect 65736 13572 65740 13628
rect 65740 13572 65796 13628
rect 65796 13572 65800 13628
rect 65736 13568 65800 13572
rect 65816 13628 65880 13632
rect 65816 13572 65820 13628
rect 65820 13572 65876 13628
rect 65876 13572 65880 13628
rect 65816 13568 65880 13572
rect 65896 13628 65960 13632
rect 65896 13572 65900 13628
rect 65900 13572 65956 13628
rect 65956 13572 65960 13628
rect 65896 13568 65960 13572
rect 19576 13084 19640 13088
rect 19576 13028 19580 13084
rect 19580 13028 19636 13084
rect 19636 13028 19640 13084
rect 19576 13024 19640 13028
rect 19656 13084 19720 13088
rect 19656 13028 19660 13084
rect 19660 13028 19716 13084
rect 19716 13028 19720 13084
rect 19656 13024 19720 13028
rect 19736 13084 19800 13088
rect 19736 13028 19740 13084
rect 19740 13028 19796 13084
rect 19796 13028 19800 13084
rect 19736 13024 19800 13028
rect 19816 13084 19880 13088
rect 19816 13028 19820 13084
rect 19820 13028 19876 13084
rect 19876 13028 19880 13084
rect 19816 13024 19880 13028
rect 50296 13084 50360 13088
rect 50296 13028 50300 13084
rect 50300 13028 50356 13084
rect 50356 13028 50360 13084
rect 50296 13024 50360 13028
rect 50376 13084 50440 13088
rect 50376 13028 50380 13084
rect 50380 13028 50436 13084
rect 50436 13028 50440 13084
rect 50376 13024 50440 13028
rect 50456 13084 50520 13088
rect 50456 13028 50460 13084
rect 50460 13028 50516 13084
rect 50516 13028 50520 13084
rect 50456 13024 50520 13028
rect 50536 13084 50600 13088
rect 50536 13028 50540 13084
rect 50540 13028 50596 13084
rect 50596 13028 50600 13084
rect 50536 13024 50600 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 65656 12540 65720 12544
rect 65656 12484 65660 12540
rect 65660 12484 65716 12540
rect 65716 12484 65720 12540
rect 65656 12480 65720 12484
rect 65736 12540 65800 12544
rect 65736 12484 65740 12540
rect 65740 12484 65796 12540
rect 65796 12484 65800 12540
rect 65736 12480 65800 12484
rect 65816 12540 65880 12544
rect 65816 12484 65820 12540
rect 65820 12484 65876 12540
rect 65876 12484 65880 12540
rect 65816 12480 65880 12484
rect 65896 12540 65960 12544
rect 65896 12484 65900 12540
rect 65900 12484 65956 12540
rect 65956 12484 65960 12540
rect 65896 12480 65960 12484
rect 19576 11996 19640 12000
rect 19576 11940 19580 11996
rect 19580 11940 19636 11996
rect 19636 11940 19640 11996
rect 19576 11936 19640 11940
rect 19656 11996 19720 12000
rect 19656 11940 19660 11996
rect 19660 11940 19716 11996
rect 19716 11940 19720 11996
rect 19656 11936 19720 11940
rect 19736 11996 19800 12000
rect 19736 11940 19740 11996
rect 19740 11940 19796 11996
rect 19796 11940 19800 11996
rect 19736 11936 19800 11940
rect 19816 11996 19880 12000
rect 19816 11940 19820 11996
rect 19820 11940 19876 11996
rect 19876 11940 19880 11996
rect 19816 11936 19880 11940
rect 50296 11996 50360 12000
rect 50296 11940 50300 11996
rect 50300 11940 50356 11996
rect 50356 11940 50360 11996
rect 50296 11936 50360 11940
rect 50376 11996 50440 12000
rect 50376 11940 50380 11996
rect 50380 11940 50436 11996
rect 50436 11940 50440 11996
rect 50376 11936 50440 11940
rect 50456 11996 50520 12000
rect 50456 11940 50460 11996
rect 50460 11940 50516 11996
rect 50516 11940 50520 11996
rect 50456 11936 50520 11940
rect 50536 11996 50600 12000
rect 50536 11940 50540 11996
rect 50540 11940 50596 11996
rect 50596 11940 50600 11996
rect 50536 11936 50600 11940
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 65656 11452 65720 11456
rect 65656 11396 65660 11452
rect 65660 11396 65716 11452
rect 65716 11396 65720 11452
rect 65656 11392 65720 11396
rect 65736 11452 65800 11456
rect 65736 11396 65740 11452
rect 65740 11396 65796 11452
rect 65796 11396 65800 11452
rect 65736 11392 65800 11396
rect 65816 11452 65880 11456
rect 65816 11396 65820 11452
rect 65820 11396 65876 11452
rect 65876 11396 65880 11452
rect 65816 11392 65880 11396
rect 65896 11452 65960 11456
rect 65896 11396 65900 11452
rect 65900 11396 65956 11452
rect 65956 11396 65960 11452
rect 65896 11392 65960 11396
rect 19576 10908 19640 10912
rect 19576 10852 19580 10908
rect 19580 10852 19636 10908
rect 19636 10852 19640 10908
rect 19576 10848 19640 10852
rect 19656 10908 19720 10912
rect 19656 10852 19660 10908
rect 19660 10852 19716 10908
rect 19716 10852 19720 10908
rect 19656 10848 19720 10852
rect 19736 10908 19800 10912
rect 19736 10852 19740 10908
rect 19740 10852 19796 10908
rect 19796 10852 19800 10908
rect 19736 10848 19800 10852
rect 19816 10908 19880 10912
rect 19816 10852 19820 10908
rect 19820 10852 19876 10908
rect 19876 10852 19880 10908
rect 19816 10848 19880 10852
rect 50296 10908 50360 10912
rect 50296 10852 50300 10908
rect 50300 10852 50356 10908
rect 50356 10852 50360 10908
rect 50296 10848 50360 10852
rect 50376 10908 50440 10912
rect 50376 10852 50380 10908
rect 50380 10852 50436 10908
rect 50436 10852 50440 10908
rect 50376 10848 50440 10852
rect 50456 10908 50520 10912
rect 50456 10852 50460 10908
rect 50460 10852 50516 10908
rect 50516 10852 50520 10908
rect 50456 10848 50520 10852
rect 50536 10908 50600 10912
rect 50536 10852 50540 10908
rect 50540 10852 50596 10908
rect 50596 10852 50600 10908
rect 50536 10848 50600 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 65656 10364 65720 10368
rect 65656 10308 65660 10364
rect 65660 10308 65716 10364
rect 65716 10308 65720 10364
rect 65656 10304 65720 10308
rect 65736 10364 65800 10368
rect 65736 10308 65740 10364
rect 65740 10308 65796 10364
rect 65796 10308 65800 10364
rect 65736 10304 65800 10308
rect 65816 10364 65880 10368
rect 65816 10308 65820 10364
rect 65820 10308 65876 10364
rect 65876 10308 65880 10364
rect 65816 10304 65880 10308
rect 65896 10364 65960 10368
rect 65896 10308 65900 10364
rect 65900 10308 65956 10364
rect 65956 10308 65960 10364
rect 65896 10304 65960 10308
rect 19576 9820 19640 9824
rect 19576 9764 19580 9820
rect 19580 9764 19636 9820
rect 19636 9764 19640 9820
rect 19576 9760 19640 9764
rect 19656 9820 19720 9824
rect 19656 9764 19660 9820
rect 19660 9764 19716 9820
rect 19716 9764 19720 9820
rect 19656 9760 19720 9764
rect 19736 9820 19800 9824
rect 19736 9764 19740 9820
rect 19740 9764 19796 9820
rect 19796 9764 19800 9820
rect 19736 9760 19800 9764
rect 19816 9820 19880 9824
rect 19816 9764 19820 9820
rect 19820 9764 19876 9820
rect 19876 9764 19880 9820
rect 19816 9760 19880 9764
rect 50296 9820 50360 9824
rect 50296 9764 50300 9820
rect 50300 9764 50356 9820
rect 50356 9764 50360 9820
rect 50296 9760 50360 9764
rect 50376 9820 50440 9824
rect 50376 9764 50380 9820
rect 50380 9764 50436 9820
rect 50436 9764 50440 9820
rect 50376 9760 50440 9764
rect 50456 9820 50520 9824
rect 50456 9764 50460 9820
rect 50460 9764 50516 9820
rect 50516 9764 50520 9820
rect 50456 9760 50520 9764
rect 50536 9820 50600 9824
rect 50536 9764 50540 9820
rect 50540 9764 50596 9820
rect 50596 9764 50600 9820
rect 50536 9760 50600 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 65656 9276 65720 9280
rect 65656 9220 65660 9276
rect 65660 9220 65716 9276
rect 65716 9220 65720 9276
rect 65656 9216 65720 9220
rect 65736 9276 65800 9280
rect 65736 9220 65740 9276
rect 65740 9220 65796 9276
rect 65796 9220 65800 9276
rect 65736 9216 65800 9220
rect 65816 9276 65880 9280
rect 65816 9220 65820 9276
rect 65820 9220 65876 9276
rect 65876 9220 65880 9276
rect 65816 9216 65880 9220
rect 65896 9276 65960 9280
rect 65896 9220 65900 9276
rect 65900 9220 65956 9276
rect 65956 9220 65960 9276
rect 65896 9216 65960 9220
rect 19576 8732 19640 8736
rect 19576 8676 19580 8732
rect 19580 8676 19636 8732
rect 19636 8676 19640 8732
rect 19576 8672 19640 8676
rect 19656 8732 19720 8736
rect 19656 8676 19660 8732
rect 19660 8676 19716 8732
rect 19716 8676 19720 8732
rect 19656 8672 19720 8676
rect 19736 8732 19800 8736
rect 19736 8676 19740 8732
rect 19740 8676 19796 8732
rect 19796 8676 19800 8732
rect 19736 8672 19800 8676
rect 19816 8732 19880 8736
rect 19816 8676 19820 8732
rect 19820 8676 19876 8732
rect 19876 8676 19880 8732
rect 19816 8672 19880 8676
rect 50296 8732 50360 8736
rect 50296 8676 50300 8732
rect 50300 8676 50356 8732
rect 50356 8676 50360 8732
rect 50296 8672 50360 8676
rect 50376 8732 50440 8736
rect 50376 8676 50380 8732
rect 50380 8676 50436 8732
rect 50436 8676 50440 8732
rect 50376 8672 50440 8676
rect 50456 8732 50520 8736
rect 50456 8676 50460 8732
rect 50460 8676 50516 8732
rect 50516 8676 50520 8732
rect 50456 8672 50520 8676
rect 50536 8732 50600 8736
rect 50536 8676 50540 8732
rect 50540 8676 50596 8732
rect 50596 8676 50600 8732
rect 50536 8672 50600 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 65656 8188 65720 8192
rect 65656 8132 65660 8188
rect 65660 8132 65716 8188
rect 65716 8132 65720 8188
rect 65656 8128 65720 8132
rect 65736 8188 65800 8192
rect 65736 8132 65740 8188
rect 65740 8132 65796 8188
rect 65796 8132 65800 8188
rect 65736 8128 65800 8132
rect 65816 8188 65880 8192
rect 65816 8132 65820 8188
rect 65820 8132 65876 8188
rect 65876 8132 65880 8188
rect 65816 8128 65880 8132
rect 65896 8188 65960 8192
rect 65896 8132 65900 8188
rect 65900 8132 65956 8188
rect 65956 8132 65960 8188
rect 65896 8128 65960 8132
rect 19576 7644 19640 7648
rect 19576 7588 19580 7644
rect 19580 7588 19636 7644
rect 19636 7588 19640 7644
rect 19576 7584 19640 7588
rect 19656 7644 19720 7648
rect 19656 7588 19660 7644
rect 19660 7588 19716 7644
rect 19716 7588 19720 7644
rect 19656 7584 19720 7588
rect 19736 7644 19800 7648
rect 19736 7588 19740 7644
rect 19740 7588 19796 7644
rect 19796 7588 19800 7644
rect 19736 7584 19800 7588
rect 19816 7644 19880 7648
rect 19816 7588 19820 7644
rect 19820 7588 19876 7644
rect 19876 7588 19880 7644
rect 19816 7584 19880 7588
rect 50296 7644 50360 7648
rect 50296 7588 50300 7644
rect 50300 7588 50356 7644
rect 50356 7588 50360 7644
rect 50296 7584 50360 7588
rect 50376 7644 50440 7648
rect 50376 7588 50380 7644
rect 50380 7588 50436 7644
rect 50436 7588 50440 7644
rect 50376 7584 50440 7588
rect 50456 7644 50520 7648
rect 50456 7588 50460 7644
rect 50460 7588 50516 7644
rect 50516 7588 50520 7644
rect 50456 7584 50520 7588
rect 50536 7644 50600 7648
rect 50536 7588 50540 7644
rect 50540 7588 50596 7644
rect 50596 7588 50600 7644
rect 50536 7584 50600 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 65656 7100 65720 7104
rect 65656 7044 65660 7100
rect 65660 7044 65716 7100
rect 65716 7044 65720 7100
rect 65656 7040 65720 7044
rect 65736 7100 65800 7104
rect 65736 7044 65740 7100
rect 65740 7044 65796 7100
rect 65796 7044 65800 7100
rect 65736 7040 65800 7044
rect 65816 7100 65880 7104
rect 65816 7044 65820 7100
rect 65820 7044 65876 7100
rect 65876 7044 65880 7100
rect 65816 7040 65880 7044
rect 65896 7100 65960 7104
rect 65896 7044 65900 7100
rect 65900 7044 65956 7100
rect 65956 7044 65960 7100
rect 65896 7040 65960 7044
rect 19576 6556 19640 6560
rect 19576 6500 19580 6556
rect 19580 6500 19636 6556
rect 19636 6500 19640 6556
rect 19576 6496 19640 6500
rect 19656 6556 19720 6560
rect 19656 6500 19660 6556
rect 19660 6500 19716 6556
rect 19716 6500 19720 6556
rect 19656 6496 19720 6500
rect 19736 6556 19800 6560
rect 19736 6500 19740 6556
rect 19740 6500 19796 6556
rect 19796 6500 19800 6556
rect 19736 6496 19800 6500
rect 19816 6556 19880 6560
rect 19816 6500 19820 6556
rect 19820 6500 19876 6556
rect 19876 6500 19880 6556
rect 19816 6496 19880 6500
rect 50296 6556 50360 6560
rect 50296 6500 50300 6556
rect 50300 6500 50356 6556
rect 50356 6500 50360 6556
rect 50296 6496 50360 6500
rect 50376 6556 50440 6560
rect 50376 6500 50380 6556
rect 50380 6500 50436 6556
rect 50436 6500 50440 6556
rect 50376 6496 50440 6500
rect 50456 6556 50520 6560
rect 50456 6500 50460 6556
rect 50460 6500 50516 6556
rect 50516 6500 50520 6556
rect 50456 6496 50520 6500
rect 50536 6556 50600 6560
rect 50536 6500 50540 6556
rect 50540 6500 50596 6556
rect 50596 6500 50600 6556
rect 50536 6496 50600 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 65656 6012 65720 6016
rect 65656 5956 65660 6012
rect 65660 5956 65716 6012
rect 65716 5956 65720 6012
rect 65656 5952 65720 5956
rect 65736 6012 65800 6016
rect 65736 5956 65740 6012
rect 65740 5956 65796 6012
rect 65796 5956 65800 6012
rect 65736 5952 65800 5956
rect 65816 6012 65880 6016
rect 65816 5956 65820 6012
rect 65820 5956 65876 6012
rect 65876 5956 65880 6012
rect 65816 5952 65880 5956
rect 65896 6012 65960 6016
rect 65896 5956 65900 6012
rect 65900 5956 65956 6012
rect 65956 5956 65960 6012
rect 65896 5952 65960 5956
rect 19576 5468 19640 5472
rect 19576 5412 19580 5468
rect 19580 5412 19636 5468
rect 19636 5412 19640 5468
rect 19576 5408 19640 5412
rect 19656 5468 19720 5472
rect 19656 5412 19660 5468
rect 19660 5412 19716 5468
rect 19716 5412 19720 5468
rect 19656 5408 19720 5412
rect 19736 5468 19800 5472
rect 19736 5412 19740 5468
rect 19740 5412 19796 5468
rect 19796 5412 19800 5468
rect 19736 5408 19800 5412
rect 19816 5468 19880 5472
rect 19816 5412 19820 5468
rect 19820 5412 19876 5468
rect 19876 5412 19880 5468
rect 19816 5408 19880 5412
rect 50296 5468 50360 5472
rect 50296 5412 50300 5468
rect 50300 5412 50356 5468
rect 50356 5412 50360 5468
rect 50296 5408 50360 5412
rect 50376 5468 50440 5472
rect 50376 5412 50380 5468
rect 50380 5412 50436 5468
rect 50436 5412 50440 5468
rect 50376 5408 50440 5412
rect 50456 5468 50520 5472
rect 50456 5412 50460 5468
rect 50460 5412 50516 5468
rect 50516 5412 50520 5468
rect 50456 5408 50520 5412
rect 50536 5468 50600 5472
rect 50536 5412 50540 5468
rect 50540 5412 50596 5468
rect 50596 5412 50600 5468
rect 50536 5408 50600 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 65656 4924 65720 4928
rect 65656 4868 65660 4924
rect 65660 4868 65716 4924
rect 65716 4868 65720 4924
rect 65656 4864 65720 4868
rect 65736 4924 65800 4928
rect 65736 4868 65740 4924
rect 65740 4868 65796 4924
rect 65796 4868 65800 4924
rect 65736 4864 65800 4868
rect 65816 4924 65880 4928
rect 65816 4868 65820 4924
rect 65820 4868 65876 4924
rect 65876 4868 65880 4924
rect 65816 4864 65880 4868
rect 65896 4924 65960 4928
rect 65896 4868 65900 4924
rect 65900 4868 65956 4924
rect 65956 4868 65960 4924
rect 65896 4864 65960 4868
rect 19576 4380 19640 4384
rect 19576 4324 19580 4380
rect 19580 4324 19636 4380
rect 19636 4324 19640 4380
rect 19576 4320 19640 4324
rect 19656 4380 19720 4384
rect 19656 4324 19660 4380
rect 19660 4324 19716 4380
rect 19716 4324 19720 4380
rect 19656 4320 19720 4324
rect 19736 4380 19800 4384
rect 19736 4324 19740 4380
rect 19740 4324 19796 4380
rect 19796 4324 19800 4380
rect 19736 4320 19800 4324
rect 19816 4380 19880 4384
rect 19816 4324 19820 4380
rect 19820 4324 19876 4380
rect 19876 4324 19880 4380
rect 19816 4320 19880 4324
rect 50296 4380 50360 4384
rect 50296 4324 50300 4380
rect 50300 4324 50356 4380
rect 50356 4324 50360 4380
rect 50296 4320 50360 4324
rect 50376 4380 50440 4384
rect 50376 4324 50380 4380
rect 50380 4324 50436 4380
rect 50436 4324 50440 4380
rect 50376 4320 50440 4324
rect 50456 4380 50520 4384
rect 50456 4324 50460 4380
rect 50460 4324 50516 4380
rect 50516 4324 50520 4380
rect 50456 4320 50520 4324
rect 50536 4380 50600 4384
rect 50536 4324 50540 4380
rect 50540 4324 50596 4380
rect 50596 4324 50600 4380
rect 50536 4320 50600 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 65656 3836 65720 3840
rect 65656 3780 65660 3836
rect 65660 3780 65716 3836
rect 65716 3780 65720 3836
rect 65656 3776 65720 3780
rect 65736 3836 65800 3840
rect 65736 3780 65740 3836
rect 65740 3780 65796 3836
rect 65796 3780 65800 3836
rect 65736 3776 65800 3780
rect 65816 3836 65880 3840
rect 65816 3780 65820 3836
rect 65820 3780 65876 3836
rect 65876 3780 65880 3836
rect 65816 3776 65880 3780
rect 65896 3836 65960 3840
rect 65896 3780 65900 3836
rect 65900 3780 65956 3836
rect 65956 3780 65960 3836
rect 65896 3776 65960 3780
rect 19576 3292 19640 3296
rect 19576 3236 19580 3292
rect 19580 3236 19636 3292
rect 19636 3236 19640 3292
rect 19576 3232 19640 3236
rect 19656 3292 19720 3296
rect 19656 3236 19660 3292
rect 19660 3236 19716 3292
rect 19716 3236 19720 3292
rect 19656 3232 19720 3236
rect 19736 3292 19800 3296
rect 19736 3236 19740 3292
rect 19740 3236 19796 3292
rect 19796 3236 19800 3292
rect 19736 3232 19800 3236
rect 19816 3292 19880 3296
rect 19816 3236 19820 3292
rect 19820 3236 19876 3292
rect 19876 3236 19880 3292
rect 19816 3232 19880 3236
rect 50296 3292 50360 3296
rect 50296 3236 50300 3292
rect 50300 3236 50356 3292
rect 50356 3236 50360 3292
rect 50296 3232 50360 3236
rect 50376 3292 50440 3296
rect 50376 3236 50380 3292
rect 50380 3236 50436 3292
rect 50436 3236 50440 3292
rect 50376 3232 50440 3236
rect 50456 3292 50520 3296
rect 50456 3236 50460 3292
rect 50460 3236 50516 3292
rect 50516 3236 50520 3292
rect 50456 3232 50520 3236
rect 50536 3292 50600 3296
rect 50536 3236 50540 3292
rect 50540 3236 50596 3292
rect 50596 3236 50600 3292
rect 50536 3232 50600 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 65656 2748 65720 2752
rect 65656 2692 65660 2748
rect 65660 2692 65716 2748
rect 65716 2692 65720 2748
rect 65656 2688 65720 2692
rect 65736 2748 65800 2752
rect 65736 2692 65740 2748
rect 65740 2692 65796 2748
rect 65796 2692 65800 2748
rect 65736 2688 65800 2692
rect 65816 2748 65880 2752
rect 65816 2692 65820 2748
rect 65820 2692 65876 2748
rect 65876 2692 65880 2748
rect 65816 2688 65880 2692
rect 65896 2748 65960 2752
rect 65896 2692 65900 2748
rect 65900 2692 65956 2748
rect 65956 2692 65960 2748
rect 65896 2688 65960 2692
rect 19576 2204 19640 2208
rect 19576 2148 19580 2204
rect 19580 2148 19636 2204
rect 19636 2148 19640 2204
rect 19576 2144 19640 2148
rect 19656 2204 19720 2208
rect 19656 2148 19660 2204
rect 19660 2148 19716 2204
rect 19716 2148 19720 2204
rect 19656 2144 19720 2148
rect 19736 2204 19800 2208
rect 19736 2148 19740 2204
rect 19740 2148 19796 2204
rect 19796 2148 19800 2204
rect 19736 2144 19800 2148
rect 19816 2204 19880 2208
rect 19816 2148 19820 2204
rect 19820 2148 19876 2204
rect 19876 2148 19880 2204
rect 19816 2144 19880 2148
rect 50296 2204 50360 2208
rect 50296 2148 50300 2204
rect 50300 2148 50356 2204
rect 50356 2148 50360 2204
rect 50296 2144 50360 2148
rect 50376 2204 50440 2208
rect 50376 2148 50380 2204
rect 50380 2148 50436 2204
rect 50436 2148 50440 2204
rect 50376 2144 50440 2148
rect 50456 2204 50520 2208
rect 50456 2148 50460 2204
rect 50460 2148 50516 2204
rect 50516 2148 50520 2204
rect 50456 2144 50520 2148
rect 50536 2204 50600 2208
rect 50536 2148 50540 2204
rect 50540 2148 50596 2204
rect 50596 2148 50600 2204
rect 50536 2144 50600 2148
<< metal4 >>
rect 4208 116992 4528 117552
rect 4208 116928 4216 116992
rect 4280 116928 4296 116992
rect 4360 116928 4376 116992
rect 4440 116928 4456 116992
rect 4520 116928 4528 116992
rect 4208 115904 4528 116928
rect 4208 115840 4216 115904
rect 4280 115840 4296 115904
rect 4360 115840 4376 115904
rect 4440 115840 4456 115904
rect 4520 115840 4528 115904
rect 4208 114816 4528 115840
rect 4208 114752 4216 114816
rect 4280 114752 4296 114816
rect 4360 114752 4376 114816
rect 4440 114752 4456 114816
rect 4520 114752 4528 114816
rect 4208 113728 4528 114752
rect 4208 113664 4216 113728
rect 4280 113664 4296 113728
rect 4360 113664 4376 113728
rect 4440 113664 4456 113728
rect 4520 113664 4528 113728
rect 4208 112640 4528 113664
rect 4208 112576 4216 112640
rect 4280 112576 4296 112640
rect 4360 112576 4376 112640
rect 4440 112576 4456 112640
rect 4520 112576 4528 112640
rect 4208 111552 4528 112576
rect 4208 111488 4216 111552
rect 4280 111488 4296 111552
rect 4360 111488 4376 111552
rect 4440 111488 4456 111552
rect 4520 111488 4528 111552
rect 4208 110464 4528 111488
rect 4208 110400 4216 110464
rect 4280 110400 4296 110464
rect 4360 110400 4376 110464
rect 4440 110400 4456 110464
rect 4520 110400 4528 110464
rect 4208 109376 4528 110400
rect 4208 109312 4216 109376
rect 4280 109312 4296 109376
rect 4360 109312 4376 109376
rect 4440 109312 4456 109376
rect 4520 109312 4528 109376
rect 4208 108288 4528 109312
rect 4208 108224 4216 108288
rect 4280 108224 4296 108288
rect 4360 108224 4376 108288
rect 4440 108224 4456 108288
rect 4520 108224 4528 108288
rect 4208 107200 4528 108224
rect 4208 107136 4216 107200
rect 4280 107136 4296 107200
rect 4360 107136 4376 107200
rect 4440 107136 4456 107200
rect 4520 107136 4528 107200
rect 4208 106112 4528 107136
rect 4208 106048 4216 106112
rect 4280 106048 4296 106112
rect 4360 106048 4376 106112
rect 4440 106048 4456 106112
rect 4520 106048 4528 106112
rect 4208 105024 4528 106048
rect 4208 104960 4216 105024
rect 4280 104960 4296 105024
rect 4360 104960 4376 105024
rect 4440 104960 4456 105024
rect 4520 104960 4528 105024
rect 4208 103936 4528 104960
rect 4208 103872 4216 103936
rect 4280 103872 4296 103936
rect 4360 103872 4376 103936
rect 4440 103872 4456 103936
rect 4520 103872 4528 103936
rect 4208 102848 4528 103872
rect 4208 102784 4216 102848
rect 4280 102784 4296 102848
rect 4360 102784 4376 102848
rect 4440 102784 4456 102848
rect 4520 102784 4528 102848
rect 4208 101760 4528 102784
rect 4208 101696 4216 101760
rect 4280 101696 4296 101760
rect 4360 101696 4376 101760
rect 4440 101696 4456 101760
rect 4520 101696 4528 101760
rect 4208 100672 4528 101696
rect 4208 100608 4216 100672
rect 4280 100608 4296 100672
rect 4360 100608 4376 100672
rect 4440 100608 4456 100672
rect 4520 100608 4528 100672
rect 4208 99584 4528 100608
rect 4208 99520 4216 99584
rect 4280 99520 4296 99584
rect 4360 99520 4376 99584
rect 4440 99520 4456 99584
rect 4520 99520 4528 99584
rect 4208 98496 4528 99520
rect 4208 98432 4216 98496
rect 4280 98432 4296 98496
rect 4360 98432 4376 98496
rect 4440 98432 4456 98496
rect 4520 98432 4528 98496
rect 4208 97484 4528 98432
rect 4208 97408 4250 97484
rect 4486 97408 4528 97484
rect 4208 97344 4216 97408
rect 4520 97344 4528 97408
rect 4208 97248 4250 97344
rect 4486 97248 4528 97344
rect 4208 96320 4528 97248
rect 4208 96256 4216 96320
rect 4280 96256 4296 96320
rect 4360 96256 4376 96320
rect 4440 96256 4456 96320
rect 4520 96256 4528 96320
rect 4208 95232 4528 96256
rect 4208 95168 4216 95232
rect 4280 95168 4296 95232
rect 4360 95168 4376 95232
rect 4440 95168 4456 95232
rect 4520 95168 4528 95232
rect 4208 94144 4528 95168
rect 4208 94080 4216 94144
rect 4280 94080 4296 94144
rect 4360 94080 4376 94144
rect 4440 94080 4456 94144
rect 4520 94080 4528 94144
rect 4208 93056 4528 94080
rect 4208 92992 4216 93056
rect 4280 92992 4296 93056
rect 4360 92992 4376 93056
rect 4440 92992 4456 93056
rect 4520 92992 4528 93056
rect 4208 91968 4528 92992
rect 4208 91904 4216 91968
rect 4280 91904 4296 91968
rect 4360 91904 4376 91968
rect 4440 91904 4456 91968
rect 4520 91904 4528 91968
rect 4208 90880 4528 91904
rect 4208 90816 4216 90880
rect 4280 90816 4296 90880
rect 4360 90816 4376 90880
rect 4440 90816 4456 90880
rect 4520 90816 4528 90880
rect 4208 89792 4528 90816
rect 4208 89728 4216 89792
rect 4280 89728 4296 89792
rect 4360 89728 4376 89792
rect 4440 89728 4456 89792
rect 4520 89728 4528 89792
rect 4208 88704 4528 89728
rect 4208 88640 4216 88704
rect 4280 88640 4296 88704
rect 4360 88640 4376 88704
rect 4440 88640 4456 88704
rect 4520 88640 4528 88704
rect 4208 87616 4528 88640
rect 4208 87552 4216 87616
rect 4280 87552 4296 87616
rect 4360 87552 4376 87616
rect 4440 87552 4456 87616
rect 4520 87552 4528 87616
rect 4208 86528 4528 87552
rect 4208 86464 4216 86528
rect 4280 86464 4296 86528
rect 4360 86464 4376 86528
rect 4440 86464 4456 86528
rect 4520 86464 4528 86528
rect 4208 85440 4528 86464
rect 4208 85376 4216 85440
rect 4280 85376 4296 85440
rect 4360 85376 4376 85440
rect 4440 85376 4456 85440
rect 4520 85376 4528 85440
rect 4208 84352 4528 85376
rect 4208 84288 4216 84352
rect 4280 84288 4296 84352
rect 4360 84288 4376 84352
rect 4440 84288 4456 84352
rect 4520 84288 4528 84352
rect 4208 83264 4528 84288
rect 4208 83200 4216 83264
rect 4280 83200 4296 83264
rect 4360 83200 4376 83264
rect 4440 83200 4456 83264
rect 4520 83200 4528 83264
rect 4208 82176 4528 83200
rect 4208 82112 4216 82176
rect 4280 82112 4296 82176
rect 4360 82112 4376 82176
rect 4440 82112 4456 82176
rect 4520 82112 4528 82176
rect 4208 81088 4528 82112
rect 4208 81024 4216 81088
rect 4280 81024 4296 81088
rect 4360 81024 4376 81088
rect 4440 81024 4456 81088
rect 4520 81024 4528 81088
rect 4208 80000 4528 81024
rect 4208 79936 4216 80000
rect 4280 79936 4296 80000
rect 4360 79936 4376 80000
rect 4440 79936 4456 80000
rect 4520 79936 4528 80000
rect 4208 78912 4528 79936
rect 4208 78848 4216 78912
rect 4280 78848 4296 78912
rect 4360 78848 4376 78912
rect 4440 78848 4456 78912
rect 4520 78848 4528 78912
rect 4208 77824 4528 78848
rect 4208 77760 4216 77824
rect 4280 77760 4296 77824
rect 4360 77760 4376 77824
rect 4440 77760 4456 77824
rect 4520 77760 4528 77824
rect 4208 76736 4528 77760
rect 4208 76672 4216 76736
rect 4280 76672 4296 76736
rect 4360 76672 4376 76736
rect 4440 76672 4456 76736
rect 4520 76672 4528 76736
rect 4208 75648 4528 76672
rect 4208 75584 4216 75648
rect 4280 75584 4296 75648
rect 4360 75584 4376 75648
rect 4440 75584 4456 75648
rect 4520 75584 4528 75648
rect 4208 74560 4528 75584
rect 4208 74496 4216 74560
rect 4280 74496 4296 74560
rect 4360 74496 4376 74560
rect 4440 74496 4456 74560
rect 4520 74496 4528 74560
rect 4208 73472 4528 74496
rect 4208 73408 4216 73472
rect 4280 73408 4296 73472
rect 4360 73408 4376 73472
rect 4440 73408 4456 73472
rect 4520 73408 4528 73472
rect 4208 72384 4528 73408
rect 4208 72320 4216 72384
rect 4280 72320 4296 72384
rect 4360 72320 4376 72384
rect 4440 72320 4456 72384
rect 4520 72320 4528 72384
rect 4208 71296 4528 72320
rect 4208 71232 4216 71296
rect 4280 71232 4296 71296
rect 4360 71232 4376 71296
rect 4440 71232 4456 71296
rect 4520 71232 4528 71296
rect 4208 70208 4528 71232
rect 4208 70144 4216 70208
rect 4280 70144 4296 70208
rect 4360 70144 4376 70208
rect 4440 70144 4456 70208
rect 4520 70144 4528 70208
rect 4208 69120 4528 70144
rect 4208 69056 4216 69120
rect 4280 69056 4296 69120
rect 4360 69056 4376 69120
rect 4440 69056 4456 69120
rect 4520 69056 4528 69120
rect 4208 68032 4528 69056
rect 4208 67968 4216 68032
rect 4280 67968 4296 68032
rect 4360 67968 4376 68032
rect 4440 67968 4456 68032
rect 4520 67968 4528 68032
rect 4208 66944 4528 67968
rect 4208 66880 4216 66944
rect 4280 66880 4296 66944
rect 4360 66880 4376 66944
rect 4440 66880 4456 66944
rect 4520 66880 4528 66944
rect 4208 66848 4528 66880
rect 4208 66612 4250 66848
rect 4486 66612 4528 66848
rect 4208 65856 4528 66612
rect 4208 65792 4216 65856
rect 4280 65792 4296 65856
rect 4360 65792 4376 65856
rect 4440 65792 4456 65856
rect 4520 65792 4528 65856
rect 4208 64768 4528 65792
rect 4208 64704 4216 64768
rect 4280 64704 4296 64768
rect 4360 64704 4376 64768
rect 4440 64704 4456 64768
rect 4520 64704 4528 64768
rect 4208 63680 4528 64704
rect 4208 63616 4216 63680
rect 4280 63616 4296 63680
rect 4360 63616 4376 63680
rect 4440 63616 4456 63680
rect 4520 63616 4528 63680
rect 4208 62592 4528 63616
rect 4208 62528 4216 62592
rect 4280 62528 4296 62592
rect 4360 62528 4376 62592
rect 4440 62528 4456 62592
rect 4520 62528 4528 62592
rect 4208 61504 4528 62528
rect 4208 61440 4216 61504
rect 4280 61440 4296 61504
rect 4360 61440 4376 61504
rect 4440 61440 4456 61504
rect 4520 61440 4528 61504
rect 4208 60416 4528 61440
rect 4208 60352 4216 60416
rect 4280 60352 4296 60416
rect 4360 60352 4376 60416
rect 4440 60352 4456 60416
rect 4520 60352 4528 60416
rect 4208 59328 4528 60352
rect 4208 59264 4216 59328
rect 4280 59264 4296 59328
rect 4360 59264 4376 59328
rect 4440 59264 4456 59328
rect 4520 59264 4528 59328
rect 4208 58240 4528 59264
rect 4208 58176 4216 58240
rect 4280 58176 4296 58240
rect 4360 58176 4376 58240
rect 4440 58176 4456 58240
rect 4520 58176 4528 58240
rect 4208 57152 4528 58176
rect 4208 57088 4216 57152
rect 4280 57088 4296 57152
rect 4360 57088 4376 57152
rect 4440 57088 4456 57152
rect 4520 57088 4528 57152
rect 4208 56064 4528 57088
rect 4208 56000 4216 56064
rect 4280 56000 4296 56064
rect 4360 56000 4376 56064
rect 4440 56000 4456 56064
rect 4520 56000 4528 56064
rect 4208 54976 4528 56000
rect 4208 54912 4216 54976
rect 4280 54912 4296 54976
rect 4360 54912 4376 54976
rect 4440 54912 4456 54976
rect 4520 54912 4528 54976
rect 4208 53888 4528 54912
rect 4208 53824 4216 53888
rect 4280 53824 4296 53888
rect 4360 53824 4376 53888
rect 4440 53824 4456 53888
rect 4520 53824 4528 53888
rect 4208 52800 4528 53824
rect 4208 52736 4216 52800
rect 4280 52736 4296 52800
rect 4360 52736 4376 52800
rect 4440 52736 4456 52800
rect 4520 52736 4528 52800
rect 4208 51712 4528 52736
rect 4208 51648 4216 51712
rect 4280 51648 4296 51712
rect 4360 51648 4376 51712
rect 4440 51648 4456 51712
rect 4520 51648 4528 51712
rect 4208 50624 4528 51648
rect 4208 50560 4216 50624
rect 4280 50560 4296 50624
rect 4360 50560 4376 50624
rect 4440 50560 4456 50624
rect 4520 50560 4528 50624
rect 4208 49536 4528 50560
rect 4208 49472 4216 49536
rect 4280 49472 4296 49536
rect 4360 49472 4376 49536
rect 4440 49472 4456 49536
rect 4520 49472 4528 49536
rect 4208 48448 4528 49472
rect 4208 48384 4216 48448
rect 4280 48384 4296 48448
rect 4360 48384 4376 48448
rect 4440 48384 4456 48448
rect 4520 48384 4528 48448
rect 4208 47360 4528 48384
rect 4208 47296 4216 47360
rect 4280 47296 4296 47360
rect 4360 47296 4376 47360
rect 4440 47296 4456 47360
rect 4520 47296 4528 47360
rect 4208 46272 4528 47296
rect 4208 46208 4216 46272
rect 4280 46208 4296 46272
rect 4360 46208 4376 46272
rect 4440 46208 4456 46272
rect 4520 46208 4528 46272
rect 4208 45184 4528 46208
rect 4208 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4528 45184
rect 4208 44096 4528 45120
rect 4208 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4528 44096
rect 4208 43008 4528 44032
rect 4208 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4528 43008
rect 4208 41920 4528 42944
rect 4208 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4528 41920
rect 4208 40832 4528 41856
rect 4208 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4528 40832
rect 4208 39744 4528 40768
rect 4208 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4528 39744
rect 4208 38656 4528 39680
rect 4208 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4528 38656
rect 4208 37568 4528 38592
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 36212 4528 36416
rect 4208 35976 4250 36212
rect 4486 35976 4528 36212
rect 4208 35392 4528 35976
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 5576 4528 5952
rect 4208 5340 4250 5576
rect 4486 5340 4528 5576
rect 4208 4928 4528 5340
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 19568 117536 19888 117552
rect 19568 117472 19576 117536
rect 19640 117472 19656 117536
rect 19720 117472 19736 117536
rect 19800 117472 19816 117536
rect 19880 117472 19888 117536
rect 19568 116448 19888 117472
rect 19568 116384 19576 116448
rect 19640 116384 19656 116448
rect 19720 116384 19736 116448
rect 19800 116384 19816 116448
rect 19880 116384 19888 116448
rect 19568 115360 19888 116384
rect 19568 115296 19576 115360
rect 19640 115296 19656 115360
rect 19720 115296 19736 115360
rect 19800 115296 19816 115360
rect 19880 115296 19888 115360
rect 19568 114272 19888 115296
rect 19568 114208 19576 114272
rect 19640 114208 19656 114272
rect 19720 114208 19736 114272
rect 19800 114208 19816 114272
rect 19880 114208 19888 114272
rect 19568 113184 19888 114208
rect 19568 113120 19576 113184
rect 19640 113120 19656 113184
rect 19720 113120 19736 113184
rect 19800 113120 19816 113184
rect 19880 113120 19888 113184
rect 19568 112802 19888 113120
rect 19568 112566 19610 112802
rect 19846 112566 19888 112802
rect 19568 112096 19888 112566
rect 19568 112032 19576 112096
rect 19640 112032 19656 112096
rect 19720 112032 19736 112096
rect 19800 112032 19816 112096
rect 19880 112032 19888 112096
rect 19568 111008 19888 112032
rect 19568 110944 19576 111008
rect 19640 110944 19656 111008
rect 19720 110944 19736 111008
rect 19800 110944 19816 111008
rect 19880 110944 19888 111008
rect 19568 109920 19888 110944
rect 19568 109856 19576 109920
rect 19640 109856 19656 109920
rect 19720 109856 19736 109920
rect 19800 109856 19816 109920
rect 19880 109856 19888 109920
rect 19568 108832 19888 109856
rect 19568 108768 19576 108832
rect 19640 108768 19656 108832
rect 19720 108768 19736 108832
rect 19800 108768 19816 108832
rect 19880 108768 19888 108832
rect 19568 107744 19888 108768
rect 19568 107680 19576 107744
rect 19640 107680 19656 107744
rect 19720 107680 19736 107744
rect 19800 107680 19816 107744
rect 19880 107680 19888 107744
rect 19568 106656 19888 107680
rect 19568 106592 19576 106656
rect 19640 106592 19656 106656
rect 19720 106592 19736 106656
rect 19800 106592 19816 106656
rect 19880 106592 19888 106656
rect 19568 105568 19888 106592
rect 19568 105504 19576 105568
rect 19640 105504 19656 105568
rect 19720 105504 19736 105568
rect 19800 105504 19816 105568
rect 19880 105504 19888 105568
rect 19568 104480 19888 105504
rect 19568 104416 19576 104480
rect 19640 104416 19656 104480
rect 19720 104416 19736 104480
rect 19800 104416 19816 104480
rect 19880 104416 19888 104480
rect 19568 103392 19888 104416
rect 19568 103328 19576 103392
rect 19640 103328 19656 103392
rect 19720 103328 19736 103392
rect 19800 103328 19816 103392
rect 19880 103328 19888 103392
rect 19568 102304 19888 103328
rect 19568 102240 19576 102304
rect 19640 102240 19656 102304
rect 19720 102240 19736 102304
rect 19800 102240 19816 102304
rect 19880 102240 19888 102304
rect 19568 101216 19888 102240
rect 19568 101152 19576 101216
rect 19640 101152 19656 101216
rect 19720 101152 19736 101216
rect 19800 101152 19816 101216
rect 19880 101152 19888 101216
rect 19568 100128 19888 101152
rect 19568 100064 19576 100128
rect 19640 100064 19656 100128
rect 19720 100064 19736 100128
rect 19800 100064 19816 100128
rect 19880 100064 19888 100128
rect 19568 99040 19888 100064
rect 19568 98976 19576 99040
rect 19640 98976 19656 99040
rect 19720 98976 19736 99040
rect 19800 98976 19816 99040
rect 19880 98976 19888 99040
rect 19568 97952 19888 98976
rect 19568 97888 19576 97952
rect 19640 97888 19656 97952
rect 19720 97888 19736 97952
rect 19800 97888 19816 97952
rect 19880 97888 19888 97952
rect 19568 96864 19888 97888
rect 19568 96800 19576 96864
rect 19640 96800 19656 96864
rect 19720 96800 19736 96864
rect 19800 96800 19816 96864
rect 19880 96800 19888 96864
rect 19568 95776 19888 96800
rect 19568 95712 19576 95776
rect 19640 95712 19656 95776
rect 19720 95712 19736 95776
rect 19800 95712 19816 95776
rect 19880 95712 19888 95776
rect 19568 94688 19888 95712
rect 19568 94624 19576 94688
rect 19640 94624 19656 94688
rect 19720 94624 19736 94688
rect 19800 94624 19816 94688
rect 19880 94624 19888 94688
rect 19568 93600 19888 94624
rect 19568 93536 19576 93600
rect 19640 93536 19656 93600
rect 19720 93536 19736 93600
rect 19800 93536 19816 93600
rect 19880 93536 19888 93600
rect 19568 92512 19888 93536
rect 19568 92448 19576 92512
rect 19640 92448 19656 92512
rect 19720 92448 19736 92512
rect 19800 92448 19816 92512
rect 19880 92448 19888 92512
rect 19568 91424 19888 92448
rect 19568 91360 19576 91424
rect 19640 91360 19656 91424
rect 19720 91360 19736 91424
rect 19800 91360 19816 91424
rect 19880 91360 19888 91424
rect 19568 90336 19888 91360
rect 19568 90272 19576 90336
rect 19640 90272 19656 90336
rect 19720 90272 19736 90336
rect 19800 90272 19816 90336
rect 19880 90272 19888 90336
rect 19568 89248 19888 90272
rect 19568 89184 19576 89248
rect 19640 89184 19656 89248
rect 19720 89184 19736 89248
rect 19800 89184 19816 89248
rect 19880 89184 19888 89248
rect 19568 88160 19888 89184
rect 19568 88096 19576 88160
rect 19640 88096 19656 88160
rect 19720 88096 19736 88160
rect 19800 88096 19816 88160
rect 19880 88096 19888 88160
rect 19568 87072 19888 88096
rect 19568 87008 19576 87072
rect 19640 87008 19656 87072
rect 19720 87008 19736 87072
rect 19800 87008 19816 87072
rect 19880 87008 19888 87072
rect 19568 85984 19888 87008
rect 19568 85920 19576 85984
rect 19640 85920 19656 85984
rect 19720 85920 19736 85984
rect 19800 85920 19816 85984
rect 19880 85920 19888 85984
rect 19568 84896 19888 85920
rect 19568 84832 19576 84896
rect 19640 84832 19656 84896
rect 19720 84832 19736 84896
rect 19800 84832 19816 84896
rect 19880 84832 19888 84896
rect 19568 83808 19888 84832
rect 19568 83744 19576 83808
rect 19640 83744 19656 83808
rect 19720 83744 19736 83808
rect 19800 83744 19816 83808
rect 19880 83744 19888 83808
rect 19568 82720 19888 83744
rect 19568 82656 19576 82720
rect 19640 82656 19656 82720
rect 19720 82656 19736 82720
rect 19800 82656 19816 82720
rect 19880 82656 19888 82720
rect 19568 82166 19888 82656
rect 19568 81930 19610 82166
rect 19846 81930 19888 82166
rect 19568 81632 19888 81930
rect 19568 81568 19576 81632
rect 19640 81568 19656 81632
rect 19720 81568 19736 81632
rect 19800 81568 19816 81632
rect 19880 81568 19888 81632
rect 19568 80544 19888 81568
rect 19568 80480 19576 80544
rect 19640 80480 19656 80544
rect 19720 80480 19736 80544
rect 19800 80480 19816 80544
rect 19880 80480 19888 80544
rect 19568 79456 19888 80480
rect 19568 79392 19576 79456
rect 19640 79392 19656 79456
rect 19720 79392 19736 79456
rect 19800 79392 19816 79456
rect 19880 79392 19888 79456
rect 19568 78368 19888 79392
rect 19568 78304 19576 78368
rect 19640 78304 19656 78368
rect 19720 78304 19736 78368
rect 19800 78304 19816 78368
rect 19880 78304 19888 78368
rect 19568 77280 19888 78304
rect 19568 77216 19576 77280
rect 19640 77216 19656 77280
rect 19720 77216 19736 77280
rect 19800 77216 19816 77280
rect 19880 77216 19888 77280
rect 19568 76192 19888 77216
rect 19568 76128 19576 76192
rect 19640 76128 19656 76192
rect 19720 76128 19736 76192
rect 19800 76128 19816 76192
rect 19880 76128 19888 76192
rect 19568 75104 19888 76128
rect 19568 75040 19576 75104
rect 19640 75040 19656 75104
rect 19720 75040 19736 75104
rect 19800 75040 19816 75104
rect 19880 75040 19888 75104
rect 19568 74016 19888 75040
rect 19568 73952 19576 74016
rect 19640 73952 19656 74016
rect 19720 73952 19736 74016
rect 19800 73952 19816 74016
rect 19880 73952 19888 74016
rect 19568 72928 19888 73952
rect 19568 72864 19576 72928
rect 19640 72864 19656 72928
rect 19720 72864 19736 72928
rect 19800 72864 19816 72928
rect 19880 72864 19888 72928
rect 19568 71840 19888 72864
rect 19568 71776 19576 71840
rect 19640 71776 19656 71840
rect 19720 71776 19736 71840
rect 19800 71776 19816 71840
rect 19880 71776 19888 71840
rect 19568 70752 19888 71776
rect 19568 70688 19576 70752
rect 19640 70688 19656 70752
rect 19720 70688 19736 70752
rect 19800 70688 19816 70752
rect 19880 70688 19888 70752
rect 19568 69664 19888 70688
rect 19568 69600 19576 69664
rect 19640 69600 19656 69664
rect 19720 69600 19736 69664
rect 19800 69600 19816 69664
rect 19880 69600 19888 69664
rect 19568 68576 19888 69600
rect 19568 68512 19576 68576
rect 19640 68512 19656 68576
rect 19720 68512 19736 68576
rect 19800 68512 19816 68576
rect 19880 68512 19888 68576
rect 19568 67488 19888 68512
rect 19568 67424 19576 67488
rect 19640 67424 19656 67488
rect 19720 67424 19736 67488
rect 19800 67424 19816 67488
rect 19880 67424 19888 67488
rect 19568 66400 19888 67424
rect 19568 66336 19576 66400
rect 19640 66336 19656 66400
rect 19720 66336 19736 66400
rect 19800 66336 19816 66400
rect 19880 66336 19888 66400
rect 19568 65312 19888 66336
rect 19568 65248 19576 65312
rect 19640 65248 19656 65312
rect 19720 65248 19736 65312
rect 19800 65248 19816 65312
rect 19880 65248 19888 65312
rect 19568 64224 19888 65248
rect 19568 64160 19576 64224
rect 19640 64160 19656 64224
rect 19720 64160 19736 64224
rect 19800 64160 19816 64224
rect 19880 64160 19888 64224
rect 19568 63136 19888 64160
rect 19568 63072 19576 63136
rect 19640 63072 19656 63136
rect 19720 63072 19736 63136
rect 19800 63072 19816 63136
rect 19880 63072 19888 63136
rect 19568 62048 19888 63072
rect 19568 61984 19576 62048
rect 19640 61984 19656 62048
rect 19720 61984 19736 62048
rect 19800 61984 19816 62048
rect 19880 61984 19888 62048
rect 19568 60960 19888 61984
rect 19568 60896 19576 60960
rect 19640 60896 19656 60960
rect 19720 60896 19736 60960
rect 19800 60896 19816 60960
rect 19880 60896 19888 60960
rect 19568 59872 19888 60896
rect 19568 59808 19576 59872
rect 19640 59808 19656 59872
rect 19720 59808 19736 59872
rect 19800 59808 19816 59872
rect 19880 59808 19888 59872
rect 19568 58784 19888 59808
rect 19568 58720 19576 58784
rect 19640 58720 19656 58784
rect 19720 58720 19736 58784
rect 19800 58720 19816 58784
rect 19880 58720 19888 58784
rect 19568 57696 19888 58720
rect 19568 57632 19576 57696
rect 19640 57632 19656 57696
rect 19720 57632 19736 57696
rect 19800 57632 19816 57696
rect 19880 57632 19888 57696
rect 19568 56608 19888 57632
rect 19568 56544 19576 56608
rect 19640 56544 19656 56608
rect 19720 56544 19736 56608
rect 19800 56544 19816 56608
rect 19880 56544 19888 56608
rect 19568 55520 19888 56544
rect 19568 55456 19576 55520
rect 19640 55456 19656 55520
rect 19720 55456 19736 55520
rect 19800 55456 19816 55520
rect 19880 55456 19888 55520
rect 19568 54432 19888 55456
rect 19568 54368 19576 54432
rect 19640 54368 19656 54432
rect 19720 54368 19736 54432
rect 19800 54368 19816 54432
rect 19880 54368 19888 54432
rect 19568 53344 19888 54368
rect 19568 53280 19576 53344
rect 19640 53280 19656 53344
rect 19720 53280 19736 53344
rect 19800 53280 19816 53344
rect 19880 53280 19888 53344
rect 19568 52256 19888 53280
rect 19568 52192 19576 52256
rect 19640 52192 19656 52256
rect 19720 52192 19736 52256
rect 19800 52192 19816 52256
rect 19880 52192 19888 52256
rect 19568 51530 19888 52192
rect 19568 51294 19610 51530
rect 19846 51294 19888 51530
rect 19568 51168 19888 51294
rect 19568 51104 19576 51168
rect 19640 51104 19656 51168
rect 19720 51104 19736 51168
rect 19800 51104 19816 51168
rect 19880 51104 19888 51168
rect 19568 50080 19888 51104
rect 19568 50016 19576 50080
rect 19640 50016 19656 50080
rect 19720 50016 19736 50080
rect 19800 50016 19816 50080
rect 19880 50016 19888 50080
rect 19568 48992 19888 50016
rect 19568 48928 19576 48992
rect 19640 48928 19656 48992
rect 19720 48928 19736 48992
rect 19800 48928 19816 48992
rect 19880 48928 19888 48992
rect 19568 47904 19888 48928
rect 19568 47840 19576 47904
rect 19640 47840 19656 47904
rect 19720 47840 19736 47904
rect 19800 47840 19816 47904
rect 19880 47840 19888 47904
rect 19568 46816 19888 47840
rect 19568 46752 19576 46816
rect 19640 46752 19656 46816
rect 19720 46752 19736 46816
rect 19800 46752 19816 46816
rect 19880 46752 19888 46816
rect 19568 45728 19888 46752
rect 19568 45664 19576 45728
rect 19640 45664 19656 45728
rect 19720 45664 19736 45728
rect 19800 45664 19816 45728
rect 19880 45664 19888 45728
rect 19568 44640 19888 45664
rect 19568 44576 19576 44640
rect 19640 44576 19656 44640
rect 19720 44576 19736 44640
rect 19800 44576 19816 44640
rect 19880 44576 19888 44640
rect 19568 43552 19888 44576
rect 19568 43488 19576 43552
rect 19640 43488 19656 43552
rect 19720 43488 19736 43552
rect 19800 43488 19816 43552
rect 19880 43488 19888 43552
rect 19568 42464 19888 43488
rect 19568 42400 19576 42464
rect 19640 42400 19656 42464
rect 19720 42400 19736 42464
rect 19800 42400 19816 42464
rect 19880 42400 19888 42464
rect 19568 41376 19888 42400
rect 19568 41312 19576 41376
rect 19640 41312 19656 41376
rect 19720 41312 19736 41376
rect 19800 41312 19816 41376
rect 19880 41312 19888 41376
rect 19568 40288 19888 41312
rect 19568 40224 19576 40288
rect 19640 40224 19656 40288
rect 19720 40224 19736 40288
rect 19800 40224 19816 40288
rect 19880 40224 19888 40288
rect 19568 39200 19888 40224
rect 19568 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19888 39200
rect 19568 38112 19888 39136
rect 19568 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19888 38112
rect 19568 37024 19888 38048
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 35936 19888 36960
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 34848 19888 35872
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 33760 19888 34784
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 32672 19888 33696
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 31584 19888 32608
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 30496 19888 31520
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 29408 19888 30432
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 28320 19888 29344
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 27232 19888 28256
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 26144 19888 27168
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 25056 19888 26080
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 23968 19888 24992
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 22880 19888 23904
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 21792 19888 22816
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 20894 19888 21728
rect 19568 20704 19610 20894
rect 19846 20704 19888 20894
rect 19568 20640 19576 20704
rect 19640 20640 19656 20658
rect 19720 20640 19736 20658
rect 19800 20640 19816 20658
rect 19880 20640 19888 20704
rect 19568 19616 19888 20640
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 18528 19888 19552
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 17440 19888 18464
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 16352 19888 17376
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 15264 19888 16288
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 14176 19888 15200
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 13088 19888 14112
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 12000 19888 13024
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 10912 19888 11936
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 9824 19888 10848
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 8736 19888 9760
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 7648 19888 8672
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 6560 19888 7584
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 5472 19888 6496
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 4384 19888 5408
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 3296 19888 4320
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19568 2208 19888 3232
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2128 19888 2144
rect 34928 116992 35248 117552
rect 34928 116928 34936 116992
rect 35000 116928 35016 116992
rect 35080 116928 35096 116992
rect 35160 116928 35176 116992
rect 35240 116928 35248 116992
rect 34928 115904 35248 116928
rect 34928 115840 34936 115904
rect 35000 115840 35016 115904
rect 35080 115840 35096 115904
rect 35160 115840 35176 115904
rect 35240 115840 35248 115904
rect 34928 114816 35248 115840
rect 34928 114752 34936 114816
rect 35000 114752 35016 114816
rect 35080 114752 35096 114816
rect 35160 114752 35176 114816
rect 35240 114752 35248 114816
rect 34928 113728 35248 114752
rect 34928 113664 34936 113728
rect 35000 113664 35016 113728
rect 35080 113664 35096 113728
rect 35160 113664 35176 113728
rect 35240 113664 35248 113728
rect 34928 112640 35248 113664
rect 34928 112576 34936 112640
rect 35000 112576 35016 112640
rect 35080 112576 35096 112640
rect 35160 112576 35176 112640
rect 35240 112576 35248 112640
rect 34928 111552 35248 112576
rect 34928 111488 34936 111552
rect 35000 111488 35016 111552
rect 35080 111488 35096 111552
rect 35160 111488 35176 111552
rect 35240 111488 35248 111552
rect 34928 110464 35248 111488
rect 34928 110400 34936 110464
rect 35000 110400 35016 110464
rect 35080 110400 35096 110464
rect 35160 110400 35176 110464
rect 35240 110400 35248 110464
rect 34928 109376 35248 110400
rect 34928 109312 34936 109376
rect 35000 109312 35016 109376
rect 35080 109312 35096 109376
rect 35160 109312 35176 109376
rect 35240 109312 35248 109376
rect 34928 108288 35248 109312
rect 34928 108224 34936 108288
rect 35000 108224 35016 108288
rect 35080 108224 35096 108288
rect 35160 108224 35176 108288
rect 35240 108224 35248 108288
rect 34928 107200 35248 108224
rect 34928 107136 34936 107200
rect 35000 107136 35016 107200
rect 35080 107136 35096 107200
rect 35160 107136 35176 107200
rect 35240 107136 35248 107200
rect 34928 106112 35248 107136
rect 34928 106048 34936 106112
rect 35000 106048 35016 106112
rect 35080 106048 35096 106112
rect 35160 106048 35176 106112
rect 35240 106048 35248 106112
rect 34928 105024 35248 106048
rect 34928 104960 34936 105024
rect 35000 104960 35016 105024
rect 35080 104960 35096 105024
rect 35160 104960 35176 105024
rect 35240 104960 35248 105024
rect 34928 103936 35248 104960
rect 34928 103872 34936 103936
rect 35000 103872 35016 103936
rect 35080 103872 35096 103936
rect 35160 103872 35176 103936
rect 35240 103872 35248 103936
rect 34928 102848 35248 103872
rect 34928 102784 34936 102848
rect 35000 102784 35016 102848
rect 35080 102784 35096 102848
rect 35160 102784 35176 102848
rect 35240 102784 35248 102848
rect 34928 101760 35248 102784
rect 34928 101696 34936 101760
rect 35000 101696 35016 101760
rect 35080 101696 35096 101760
rect 35160 101696 35176 101760
rect 35240 101696 35248 101760
rect 34928 100672 35248 101696
rect 34928 100608 34936 100672
rect 35000 100608 35016 100672
rect 35080 100608 35096 100672
rect 35160 100608 35176 100672
rect 35240 100608 35248 100672
rect 34928 99584 35248 100608
rect 34928 99520 34936 99584
rect 35000 99520 35016 99584
rect 35080 99520 35096 99584
rect 35160 99520 35176 99584
rect 35240 99520 35248 99584
rect 34928 98496 35248 99520
rect 34928 98432 34936 98496
rect 35000 98432 35016 98496
rect 35080 98432 35096 98496
rect 35160 98432 35176 98496
rect 35240 98432 35248 98496
rect 34928 97484 35248 98432
rect 34928 97408 34970 97484
rect 35206 97408 35248 97484
rect 34928 97344 34936 97408
rect 35240 97344 35248 97408
rect 34928 97248 34970 97344
rect 35206 97248 35248 97344
rect 34928 96320 35248 97248
rect 34928 96256 34936 96320
rect 35000 96256 35016 96320
rect 35080 96256 35096 96320
rect 35160 96256 35176 96320
rect 35240 96256 35248 96320
rect 34928 95232 35248 96256
rect 34928 95168 34936 95232
rect 35000 95168 35016 95232
rect 35080 95168 35096 95232
rect 35160 95168 35176 95232
rect 35240 95168 35248 95232
rect 34928 94144 35248 95168
rect 34928 94080 34936 94144
rect 35000 94080 35016 94144
rect 35080 94080 35096 94144
rect 35160 94080 35176 94144
rect 35240 94080 35248 94144
rect 34928 93056 35248 94080
rect 34928 92992 34936 93056
rect 35000 92992 35016 93056
rect 35080 92992 35096 93056
rect 35160 92992 35176 93056
rect 35240 92992 35248 93056
rect 34928 91968 35248 92992
rect 34928 91904 34936 91968
rect 35000 91904 35016 91968
rect 35080 91904 35096 91968
rect 35160 91904 35176 91968
rect 35240 91904 35248 91968
rect 34928 90880 35248 91904
rect 34928 90816 34936 90880
rect 35000 90816 35016 90880
rect 35080 90816 35096 90880
rect 35160 90816 35176 90880
rect 35240 90816 35248 90880
rect 34928 89792 35248 90816
rect 34928 89728 34936 89792
rect 35000 89728 35016 89792
rect 35080 89728 35096 89792
rect 35160 89728 35176 89792
rect 35240 89728 35248 89792
rect 34928 88704 35248 89728
rect 34928 88640 34936 88704
rect 35000 88640 35016 88704
rect 35080 88640 35096 88704
rect 35160 88640 35176 88704
rect 35240 88640 35248 88704
rect 34928 87616 35248 88640
rect 34928 87552 34936 87616
rect 35000 87552 35016 87616
rect 35080 87552 35096 87616
rect 35160 87552 35176 87616
rect 35240 87552 35248 87616
rect 34928 86528 35248 87552
rect 34928 86464 34936 86528
rect 35000 86464 35016 86528
rect 35080 86464 35096 86528
rect 35160 86464 35176 86528
rect 35240 86464 35248 86528
rect 34928 85440 35248 86464
rect 34928 85376 34936 85440
rect 35000 85376 35016 85440
rect 35080 85376 35096 85440
rect 35160 85376 35176 85440
rect 35240 85376 35248 85440
rect 34928 84352 35248 85376
rect 34928 84288 34936 84352
rect 35000 84288 35016 84352
rect 35080 84288 35096 84352
rect 35160 84288 35176 84352
rect 35240 84288 35248 84352
rect 34928 83264 35248 84288
rect 34928 83200 34936 83264
rect 35000 83200 35016 83264
rect 35080 83200 35096 83264
rect 35160 83200 35176 83264
rect 35240 83200 35248 83264
rect 34928 82176 35248 83200
rect 34928 82112 34936 82176
rect 35000 82112 35016 82176
rect 35080 82112 35096 82176
rect 35160 82112 35176 82176
rect 35240 82112 35248 82176
rect 34928 81088 35248 82112
rect 34928 81024 34936 81088
rect 35000 81024 35016 81088
rect 35080 81024 35096 81088
rect 35160 81024 35176 81088
rect 35240 81024 35248 81088
rect 34928 80000 35248 81024
rect 34928 79936 34936 80000
rect 35000 79936 35016 80000
rect 35080 79936 35096 80000
rect 35160 79936 35176 80000
rect 35240 79936 35248 80000
rect 34928 78912 35248 79936
rect 34928 78848 34936 78912
rect 35000 78848 35016 78912
rect 35080 78848 35096 78912
rect 35160 78848 35176 78912
rect 35240 78848 35248 78912
rect 34928 77824 35248 78848
rect 34928 77760 34936 77824
rect 35000 77760 35016 77824
rect 35080 77760 35096 77824
rect 35160 77760 35176 77824
rect 35240 77760 35248 77824
rect 34928 76736 35248 77760
rect 34928 76672 34936 76736
rect 35000 76672 35016 76736
rect 35080 76672 35096 76736
rect 35160 76672 35176 76736
rect 35240 76672 35248 76736
rect 34928 75648 35248 76672
rect 34928 75584 34936 75648
rect 35000 75584 35016 75648
rect 35080 75584 35096 75648
rect 35160 75584 35176 75648
rect 35240 75584 35248 75648
rect 34928 74560 35248 75584
rect 34928 74496 34936 74560
rect 35000 74496 35016 74560
rect 35080 74496 35096 74560
rect 35160 74496 35176 74560
rect 35240 74496 35248 74560
rect 34928 73472 35248 74496
rect 34928 73408 34936 73472
rect 35000 73408 35016 73472
rect 35080 73408 35096 73472
rect 35160 73408 35176 73472
rect 35240 73408 35248 73472
rect 34928 72384 35248 73408
rect 34928 72320 34936 72384
rect 35000 72320 35016 72384
rect 35080 72320 35096 72384
rect 35160 72320 35176 72384
rect 35240 72320 35248 72384
rect 34928 71296 35248 72320
rect 34928 71232 34936 71296
rect 35000 71232 35016 71296
rect 35080 71232 35096 71296
rect 35160 71232 35176 71296
rect 35240 71232 35248 71296
rect 34928 70208 35248 71232
rect 34928 70144 34936 70208
rect 35000 70144 35016 70208
rect 35080 70144 35096 70208
rect 35160 70144 35176 70208
rect 35240 70144 35248 70208
rect 34928 69120 35248 70144
rect 34928 69056 34936 69120
rect 35000 69056 35016 69120
rect 35080 69056 35096 69120
rect 35160 69056 35176 69120
rect 35240 69056 35248 69120
rect 34928 68032 35248 69056
rect 34928 67968 34936 68032
rect 35000 67968 35016 68032
rect 35080 67968 35096 68032
rect 35160 67968 35176 68032
rect 35240 67968 35248 68032
rect 34928 66944 35248 67968
rect 34928 66880 34936 66944
rect 35000 66880 35016 66944
rect 35080 66880 35096 66944
rect 35160 66880 35176 66944
rect 35240 66880 35248 66944
rect 34928 66848 35248 66880
rect 34928 66612 34970 66848
rect 35206 66612 35248 66848
rect 34928 65856 35248 66612
rect 34928 65792 34936 65856
rect 35000 65792 35016 65856
rect 35080 65792 35096 65856
rect 35160 65792 35176 65856
rect 35240 65792 35248 65856
rect 34928 64768 35248 65792
rect 34928 64704 34936 64768
rect 35000 64704 35016 64768
rect 35080 64704 35096 64768
rect 35160 64704 35176 64768
rect 35240 64704 35248 64768
rect 34928 63680 35248 64704
rect 34928 63616 34936 63680
rect 35000 63616 35016 63680
rect 35080 63616 35096 63680
rect 35160 63616 35176 63680
rect 35240 63616 35248 63680
rect 34928 62592 35248 63616
rect 34928 62528 34936 62592
rect 35000 62528 35016 62592
rect 35080 62528 35096 62592
rect 35160 62528 35176 62592
rect 35240 62528 35248 62592
rect 34928 61504 35248 62528
rect 34928 61440 34936 61504
rect 35000 61440 35016 61504
rect 35080 61440 35096 61504
rect 35160 61440 35176 61504
rect 35240 61440 35248 61504
rect 34928 60416 35248 61440
rect 34928 60352 34936 60416
rect 35000 60352 35016 60416
rect 35080 60352 35096 60416
rect 35160 60352 35176 60416
rect 35240 60352 35248 60416
rect 34928 59328 35248 60352
rect 34928 59264 34936 59328
rect 35000 59264 35016 59328
rect 35080 59264 35096 59328
rect 35160 59264 35176 59328
rect 35240 59264 35248 59328
rect 34928 58240 35248 59264
rect 34928 58176 34936 58240
rect 35000 58176 35016 58240
rect 35080 58176 35096 58240
rect 35160 58176 35176 58240
rect 35240 58176 35248 58240
rect 34928 57152 35248 58176
rect 34928 57088 34936 57152
rect 35000 57088 35016 57152
rect 35080 57088 35096 57152
rect 35160 57088 35176 57152
rect 35240 57088 35248 57152
rect 34928 56064 35248 57088
rect 34928 56000 34936 56064
rect 35000 56000 35016 56064
rect 35080 56000 35096 56064
rect 35160 56000 35176 56064
rect 35240 56000 35248 56064
rect 34928 54976 35248 56000
rect 34928 54912 34936 54976
rect 35000 54912 35016 54976
rect 35080 54912 35096 54976
rect 35160 54912 35176 54976
rect 35240 54912 35248 54976
rect 34928 53888 35248 54912
rect 34928 53824 34936 53888
rect 35000 53824 35016 53888
rect 35080 53824 35096 53888
rect 35160 53824 35176 53888
rect 35240 53824 35248 53888
rect 34928 52800 35248 53824
rect 34928 52736 34936 52800
rect 35000 52736 35016 52800
rect 35080 52736 35096 52800
rect 35160 52736 35176 52800
rect 35240 52736 35248 52800
rect 34928 51712 35248 52736
rect 34928 51648 34936 51712
rect 35000 51648 35016 51712
rect 35080 51648 35096 51712
rect 35160 51648 35176 51712
rect 35240 51648 35248 51712
rect 34928 50624 35248 51648
rect 34928 50560 34936 50624
rect 35000 50560 35016 50624
rect 35080 50560 35096 50624
rect 35160 50560 35176 50624
rect 35240 50560 35248 50624
rect 34928 49536 35248 50560
rect 34928 49472 34936 49536
rect 35000 49472 35016 49536
rect 35080 49472 35096 49536
rect 35160 49472 35176 49536
rect 35240 49472 35248 49536
rect 34928 48448 35248 49472
rect 34928 48384 34936 48448
rect 35000 48384 35016 48448
rect 35080 48384 35096 48448
rect 35160 48384 35176 48448
rect 35240 48384 35248 48448
rect 34928 47360 35248 48384
rect 34928 47296 34936 47360
rect 35000 47296 35016 47360
rect 35080 47296 35096 47360
rect 35160 47296 35176 47360
rect 35240 47296 35248 47360
rect 34928 46272 35248 47296
rect 34928 46208 34936 46272
rect 35000 46208 35016 46272
rect 35080 46208 35096 46272
rect 35160 46208 35176 46272
rect 35240 46208 35248 46272
rect 34928 45184 35248 46208
rect 34928 45120 34936 45184
rect 35000 45120 35016 45184
rect 35080 45120 35096 45184
rect 35160 45120 35176 45184
rect 35240 45120 35248 45184
rect 34928 44096 35248 45120
rect 34928 44032 34936 44096
rect 35000 44032 35016 44096
rect 35080 44032 35096 44096
rect 35160 44032 35176 44096
rect 35240 44032 35248 44096
rect 34928 43008 35248 44032
rect 34928 42944 34936 43008
rect 35000 42944 35016 43008
rect 35080 42944 35096 43008
rect 35160 42944 35176 43008
rect 35240 42944 35248 43008
rect 34928 41920 35248 42944
rect 34928 41856 34936 41920
rect 35000 41856 35016 41920
rect 35080 41856 35096 41920
rect 35160 41856 35176 41920
rect 35240 41856 35248 41920
rect 34928 40832 35248 41856
rect 34928 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35248 40832
rect 34928 39744 35248 40768
rect 34928 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35248 39744
rect 34928 38656 35248 39680
rect 34928 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35248 38656
rect 34928 37568 35248 38592
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 36480 35248 37504
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 36212 35248 36416
rect 34928 35976 34970 36212
rect 35206 35976 35248 36212
rect 34928 35392 35248 35976
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 34304 35248 35328
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 32128 35248 33152
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 31040 35248 32064
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 29952 35248 30976
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 28864 35248 29888
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 27776 35248 28800
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 26688 35248 27712
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 25600 35248 26624
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 24512 35248 25536
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 23424 35248 24448
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 22336 35248 23360
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 21248 35248 22272
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 20160 35248 21184
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 19072 35248 20096
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 17984 35248 19008
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 16896 35248 17920
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 14720 35248 15744
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 13632 35248 14656
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 12544 35248 13568
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 11456 35248 12480
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 9280 35248 10304
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 8192 35248 9216
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 5576 35248 5952
rect 34928 5340 34970 5576
rect 35206 5340 35248 5576
rect 34928 4928 35248 5340
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2128 35248 2688
rect 50288 117536 50608 117552
rect 50288 117472 50296 117536
rect 50360 117472 50376 117536
rect 50440 117472 50456 117536
rect 50520 117472 50536 117536
rect 50600 117472 50608 117536
rect 50288 116448 50608 117472
rect 50288 116384 50296 116448
rect 50360 116384 50376 116448
rect 50440 116384 50456 116448
rect 50520 116384 50536 116448
rect 50600 116384 50608 116448
rect 50288 115360 50608 116384
rect 50288 115296 50296 115360
rect 50360 115296 50376 115360
rect 50440 115296 50456 115360
rect 50520 115296 50536 115360
rect 50600 115296 50608 115360
rect 50288 114272 50608 115296
rect 50288 114208 50296 114272
rect 50360 114208 50376 114272
rect 50440 114208 50456 114272
rect 50520 114208 50536 114272
rect 50600 114208 50608 114272
rect 50288 113184 50608 114208
rect 50288 113120 50296 113184
rect 50360 113120 50376 113184
rect 50440 113120 50456 113184
rect 50520 113120 50536 113184
rect 50600 113120 50608 113184
rect 50288 112802 50608 113120
rect 50288 112566 50330 112802
rect 50566 112566 50608 112802
rect 50288 112096 50608 112566
rect 50288 112032 50296 112096
rect 50360 112032 50376 112096
rect 50440 112032 50456 112096
rect 50520 112032 50536 112096
rect 50600 112032 50608 112096
rect 50288 111008 50608 112032
rect 50288 110944 50296 111008
rect 50360 110944 50376 111008
rect 50440 110944 50456 111008
rect 50520 110944 50536 111008
rect 50600 110944 50608 111008
rect 50288 109920 50608 110944
rect 50288 109856 50296 109920
rect 50360 109856 50376 109920
rect 50440 109856 50456 109920
rect 50520 109856 50536 109920
rect 50600 109856 50608 109920
rect 50288 108832 50608 109856
rect 50288 108768 50296 108832
rect 50360 108768 50376 108832
rect 50440 108768 50456 108832
rect 50520 108768 50536 108832
rect 50600 108768 50608 108832
rect 50288 107744 50608 108768
rect 50288 107680 50296 107744
rect 50360 107680 50376 107744
rect 50440 107680 50456 107744
rect 50520 107680 50536 107744
rect 50600 107680 50608 107744
rect 50288 106656 50608 107680
rect 50288 106592 50296 106656
rect 50360 106592 50376 106656
rect 50440 106592 50456 106656
rect 50520 106592 50536 106656
rect 50600 106592 50608 106656
rect 50288 105568 50608 106592
rect 50288 105504 50296 105568
rect 50360 105504 50376 105568
rect 50440 105504 50456 105568
rect 50520 105504 50536 105568
rect 50600 105504 50608 105568
rect 50288 104480 50608 105504
rect 50288 104416 50296 104480
rect 50360 104416 50376 104480
rect 50440 104416 50456 104480
rect 50520 104416 50536 104480
rect 50600 104416 50608 104480
rect 50288 103392 50608 104416
rect 50288 103328 50296 103392
rect 50360 103328 50376 103392
rect 50440 103328 50456 103392
rect 50520 103328 50536 103392
rect 50600 103328 50608 103392
rect 50288 102304 50608 103328
rect 50288 102240 50296 102304
rect 50360 102240 50376 102304
rect 50440 102240 50456 102304
rect 50520 102240 50536 102304
rect 50600 102240 50608 102304
rect 50288 101216 50608 102240
rect 50288 101152 50296 101216
rect 50360 101152 50376 101216
rect 50440 101152 50456 101216
rect 50520 101152 50536 101216
rect 50600 101152 50608 101216
rect 50288 100128 50608 101152
rect 50288 100064 50296 100128
rect 50360 100064 50376 100128
rect 50440 100064 50456 100128
rect 50520 100064 50536 100128
rect 50600 100064 50608 100128
rect 50288 99040 50608 100064
rect 50288 98976 50296 99040
rect 50360 98976 50376 99040
rect 50440 98976 50456 99040
rect 50520 98976 50536 99040
rect 50600 98976 50608 99040
rect 50288 97952 50608 98976
rect 50288 97888 50296 97952
rect 50360 97888 50376 97952
rect 50440 97888 50456 97952
rect 50520 97888 50536 97952
rect 50600 97888 50608 97952
rect 50288 96864 50608 97888
rect 50288 96800 50296 96864
rect 50360 96800 50376 96864
rect 50440 96800 50456 96864
rect 50520 96800 50536 96864
rect 50600 96800 50608 96864
rect 50288 95776 50608 96800
rect 50288 95712 50296 95776
rect 50360 95712 50376 95776
rect 50440 95712 50456 95776
rect 50520 95712 50536 95776
rect 50600 95712 50608 95776
rect 50288 94688 50608 95712
rect 50288 94624 50296 94688
rect 50360 94624 50376 94688
rect 50440 94624 50456 94688
rect 50520 94624 50536 94688
rect 50600 94624 50608 94688
rect 50288 93600 50608 94624
rect 50288 93536 50296 93600
rect 50360 93536 50376 93600
rect 50440 93536 50456 93600
rect 50520 93536 50536 93600
rect 50600 93536 50608 93600
rect 50288 92512 50608 93536
rect 50288 92448 50296 92512
rect 50360 92448 50376 92512
rect 50440 92448 50456 92512
rect 50520 92448 50536 92512
rect 50600 92448 50608 92512
rect 50288 91424 50608 92448
rect 50288 91360 50296 91424
rect 50360 91360 50376 91424
rect 50440 91360 50456 91424
rect 50520 91360 50536 91424
rect 50600 91360 50608 91424
rect 50288 90336 50608 91360
rect 50288 90272 50296 90336
rect 50360 90272 50376 90336
rect 50440 90272 50456 90336
rect 50520 90272 50536 90336
rect 50600 90272 50608 90336
rect 50288 89248 50608 90272
rect 50288 89184 50296 89248
rect 50360 89184 50376 89248
rect 50440 89184 50456 89248
rect 50520 89184 50536 89248
rect 50600 89184 50608 89248
rect 50288 88160 50608 89184
rect 50288 88096 50296 88160
rect 50360 88096 50376 88160
rect 50440 88096 50456 88160
rect 50520 88096 50536 88160
rect 50600 88096 50608 88160
rect 50288 87072 50608 88096
rect 50288 87008 50296 87072
rect 50360 87008 50376 87072
rect 50440 87008 50456 87072
rect 50520 87008 50536 87072
rect 50600 87008 50608 87072
rect 50288 85984 50608 87008
rect 50288 85920 50296 85984
rect 50360 85920 50376 85984
rect 50440 85920 50456 85984
rect 50520 85920 50536 85984
rect 50600 85920 50608 85984
rect 50288 84896 50608 85920
rect 50288 84832 50296 84896
rect 50360 84832 50376 84896
rect 50440 84832 50456 84896
rect 50520 84832 50536 84896
rect 50600 84832 50608 84896
rect 50288 83808 50608 84832
rect 50288 83744 50296 83808
rect 50360 83744 50376 83808
rect 50440 83744 50456 83808
rect 50520 83744 50536 83808
rect 50600 83744 50608 83808
rect 50288 82720 50608 83744
rect 50288 82656 50296 82720
rect 50360 82656 50376 82720
rect 50440 82656 50456 82720
rect 50520 82656 50536 82720
rect 50600 82656 50608 82720
rect 50288 82166 50608 82656
rect 50288 81930 50330 82166
rect 50566 81930 50608 82166
rect 50288 81632 50608 81930
rect 50288 81568 50296 81632
rect 50360 81568 50376 81632
rect 50440 81568 50456 81632
rect 50520 81568 50536 81632
rect 50600 81568 50608 81632
rect 50288 80544 50608 81568
rect 50288 80480 50296 80544
rect 50360 80480 50376 80544
rect 50440 80480 50456 80544
rect 50520 80480 50536 80544
rect 50600 80480 50608 80544
rect 50288 79456 50608 80480
rect 50288 79392 50296 79456
rect 50360 79392 50376 79456
rect 50440 79392 50456 79456
rect 50520 79392 50536 79456
rect 50600 79392 50608 79456
rect 50288 78368 50608 79392
rect 50288 78304 50296 78368
rect 50360 78304 50376 78368
rect 50440 78304 50456 78368
rect 50520 78304 50536 78368
rect 50600 78304 50608 78368
rect 50288 77280 50608 78304
rect 50288 77216 50296 77280
rect 50360 77216 50376 77280
rect 50440 77216 50456 77280
rect 50520 77216 50536 77280
rect 50600 77216 50608 77280
rect 50288 76192 50608 77216
rect 50288 76128 50296 76192
rect 50360 76128 50376 76192
rect 50440 76128 50456 76192
rect 50520 76128 50536 76192
rect 50600 76128 50608 76192
rect 50288 75104 50608 76128
rect 50288 75040 50296 75104
rect 50360 75040 50376 75104
rect 50440 75040 50456 75104
rect 50520 75040 50536 75104
rect 50600 75040 50608 75104
rect 50288 74016 50608 75040
rect 50288 73952 50296 74016
rect 50360 73952 50376 74016
rect 50440 73952 50456 74016
rect 50520 73952 50536 74016
rect 50600 73952 50608 74016
rect 50288 72928 50608 73952
rect 50288 72864 50296 72928
rect 50360 72864 50376 72928
rect 50440 72864 50456 72928
rect 50520 72864 50536 72928
rect 50600 72864 50608 72928
rect 50288 71840 50608 72864
rect 50288 71776 50296 71840
rect 50360 71776 50376 71840
rect 50440 71776 50456 71840
rect 50520 71776 50536 71840
rect 50600 71776 50608 71840
rect 50288 70752 50608 71776
rect 50288 70688 50296 70752
rect 50360 70688 50376 70752
rect 50440 70688 50456 70752
rect 50520 70688 50536 70752
rect 50600 70688 50608 70752
rect 50288 69664 50608 70688
rect 50288 69600 50296 69664
rect 50360 69600 50376 69664
rect 50440 69600 50456 69664
rect 50520 69600 50536 69664
rect 50600 69600 50608 69664
rect 50288 68576 50608 69600
rect 50288 68512 50296 68576
rect 50360 68512 50376 68576
rect 50440 68512 50456 68576
rect 50520 68512 50536 68576
rect 50600 68512 50608 68576
rect 50288 67488 50608 68512
rect 50288 67424 50296 67488
rect 50360 67424 50376 67488
rect 50440 67424 50456 67488
rect 50520 67424 50536 67488
rect 50600 67424 50608 67488
rect 50288 66400 50608 67424
rect 50288 66336 50296 66400
rect 50360 66336 50376 66400
rect 50440 66336 50456 66400
rect 50520 66336 50536 66400
rect 50600 66336 50608 66400
rect 50288 65312 50608 66336
rect 50288 65248 50296 65312
rect 50360 65248 50376 65312
rect 50440 65248 50456 65312
rect 50520 65248 50536 65312
rect 50600 65248 50608 65312
rect 50288 64224 50608 65248
rect 50288 64160 50296 64224
rect 50360 64160 50376 64224
rect 50440 64160 50456 64224
rect 50520 64160 50536 64224
rect 50600 64160 50608 64224
rect 50288 63136 50608 64160
rect 50288 63072 50296 63136
rect 50360 63072 50376 63136
rect 50440 63072 50456 63136
rect 50520 63072 50536 63136
rect 50600 63072 50608 63136
rect 50288 62048 50608 63072
rect 50288 61984 50296 62048
rect 50360 61984 50376 62048
rect 50440 61984 50456 62048
rect 50520 61984 50536 62048
rect 50600 61984 50608 62048
rect 50288 60960 50608 61984
rect 50288 60896 50296 60960
rect 50360 60896 50376 60960
rect 50440 60896 50456 60960
rect 50520 60896 50536 60960
rect 50600 60896 50608 60960
rect 50288 59872 50608 60896
rect 50288 59808 50296 59872
rect 50360 59808 50376 59872
rect 50440 59808 50456 59872
rect 50520 59808 50536 59872
rect 50600 59808 50608 59872
rect 50288 58784 50608 59808
rect 50288 58720 50296 58784
rect 50360 58720 50376 58784
rect 50440 58720 50456 58784
rect 50520 58720 50536 58784
rect 50600 58720 50608 58784
rect 50288 57696 50608 58720
rect 50288 57632 50296 57696
rect 50360 57632 50376 57696
rect 50440 57632 50456 57696
rect 50520 57632 50536 57696
rect 50600 57632 50608 57696
rect 50288 56608 50608 57632
rect 50288 56544 50296 56608
rect 50360 56544 50376 56608
rect 50440 56544 50456 56608
rect 50520 56544 50536 56608
rect 50600 56544 50608 56608
rect 50288 55520 50608 56544
rect 50288 55456 50296 55520
rect 50360 55456 50376 55520
rect 50440 55456 50456 55520
rect 50520 55456 50536 55520
rect 50600 55456 50608 55520
rect 50288 54432 50608 55456
rect 50288 54368 50296 54432
rect 50360 54368 50376 54432
rect 50440 54368 50456 54432
rect 50520 54368 50536 54432
rect 50600 54368 50608 54432
rect 50288 53344 50608 54368
rect 50288 53280 50296 53344
rect 50360 53280 50376 53344
rect 50440 53280 50456 53344
rect 50520 53280 50536 53344
rect 50600 53280 50608 53344
rect 50288 52256 50608 53280
rect 50288 52192 50296 52256
rect 50360 52192 50376 52256
rect 50440 52192 50456 52256
rect 50520 52192 50536 52256
rect 50600 52192 50608 52256
rect 50288 51530 50608 52192
rect 50288 51294 50330 51530
rect 50566 51294 50608 51530
rect 50288 51168 50608 51294
rect 50288 51104 50296 51168
rect 50360 51104 50376 51168
rect 50440 51104 50456 51168
rect 50520 51104 50536 51168
rect 50600 51104 50608 51168
rect 50288 50080 50608 51104
rect 50288 50016 50296 50080
rect 50360 50016 50376 50080
rect 50440 50016 50456 50080
rect 50520 50016 50536 50080
rect 50600 50016 50608 50080
rect 50288 48992 50608 50016
rect 50288 48928 50296 48992
rect 50360 48928 50376 48992
rect 50440 48928 50456 48992
rect 50520 48928 50536 48992
rect 50600 48928 50608 48992
rect 50288 47904 50608 48928
rect 50288 47840 50296 47904
rect 50360 47840 50376 47904
rect 50440 47840 50456 47904
rect 50520 47840 50536 47904
rect 50600 47840 50608 47904
rect 50288 46816 50608 47840
rect 50288 46752 50296 46816
rect 50360 46752 50376 46816
rect 50440 46752 50456 46816
rect 50520 46752 50536 46816
rect 50600 46752 50608 46816
rect 50288 45728 50608 46752
rect 50288 45664 50296 45728
rect 50360 45664 50376 45728
rect 50440 45664 50456 45728
rect 50520 45664 50536 45728
rect 50600 45664 50608 45728
rect 50288 44640 50608 45664
rect 50288 44576 50296 44640
rect 50360 44576 50376 44640
rect 50440 44576 50456 44640
rect 50520 44576 50536 44640
rect 50600 44576 50608 44640
rect 50288 43552 50608 44576
rect 50288 43488 50296 43552
rect 50360 43488 50376 43552
rect 50440 43488 50456 43552
rect 50520 43488 50536 43552
rect 50600 43488 50608 43552
rect 50288 42464 50608 43488
rect 50288 42400 50296 42464
rect 50360 42400 50376 42464
rect 50440 42400 50456 42464
rect 50520 42400 50536 42464
rect 50600 42400 50608 42464
rect 50288 41376 50608 42400
rect 50288 41312 50296 41376
rect 50360 41312 50376 41376
rect 50440 41312 50456 41376
rect 50520 41312 50536 41376
rect 50600 41312 50608 41376
rect 50288 40288 50608 41312
rect 50288 40224 50296 40288
rect 50360 40224 50376 40288
rect 50440 40224 50456 40288
rect 50520 40224 50536 40288
rect 50600 40224 50608 40288
rect 50288 39200 50608 40224
rect 50288 39136 50296 39200
rect 50360 39136 50376 39200
rect 50440 39136 50456 39200
rect 50520 39136 50536 39200
rect 50600 39136 50608 39200
rect 50288 38112 50608 39136
rect 50288 38048 50296 38112
rect 50360 38048 50376 38112
rect 50440 38048 50456 38112
rect 50520 38048 50536 38112
rect 50600 38048 50608 38112
rect 50288 37024 50608 38048
rect 50288 36960 50296 37024
rect 50360 36960 50376 37024
rect 50440 36960 50456 37024
rect 50520 36960 50536 37024
rect 50600 36960 50608 37024
rect 50288 35936 50608 36960
rect 50288 35872 50296 35936
rect 50360 35872 50376 35936
rect 50440 35872 50456 35936
rect 50520 35872 50536 35936
rect 50600 35872 50608 35936
rect 50288 34848 50608 35872
rect 50288 34784 50296 34848
rect 50360 34784 50376 34848
rect 50440 34784 50456 34848
rect 50520 34784 50536 34848
rect 50600 34784 50608 34848
rect 50288 33760 50608 34784
rect 50288 33696 50296 33760
rect 50360 33696 50376 33760
rect 50440 33696 50456 33760
rect 50520 33696 50536 33760
rect 50600 33696 50608 33760
rect 50288 32672 50608 33696
rect 50288 32608 50296 32672
rect 50360 32608 50376 32672
rect 50440 32608 50456 32672
rect 50520 32608 50536 32672
rect 50600 32608 50608 32672
rect 50288 31584 50608 32608
rect 50288 31520 50296 31584
rect 50360 31520 50376 31584
rect 50440 31520 50456 31584
rect 50520 31520 50536 31584
rect 50600 31520 50608 31584
rect 50288 30496 50608 31520
rect 50288 30432 50296 30496
rect 50360 30432 50376 30496
rect 50440 30432 50456 30496
rect 50520 30432 50536 30496
rect 50600 30432 50608 30496
rect 50288 29408 50608 30432
rect 50288 29344 50296 29408
rect 50360 29344 50376 29408
rect 50440 29344 50456 29408
rect 50520 29344 50536 29408
rect 50600 29344 50608 29408
rect 50288 28320 50608 29344
rect 50288 28256 50296 28320
rect 50360 28256 50376 28320
rect 50440 28256 50456 28320
rect 50520 28256 50536 28320
rect 50600 28256 50608 28320
rect 50288 27232 50608 28256
rect 50288 27168 50296 27232
rect 50360 27168 50376 27232
rect 50440 27168 50456 27232
rect 50520 27168 50536 27232
rect 50600 27168 50608 27232
rect 50288 26144 50608 27168
rect 50288 26080 50296 26144
rect 50360 26080 50376 26144
rect 50440 26080 50456 26144
rect 50520 26080 50536 26144
rect 50600 26080 50608 26144
rect 50288 25056 50608 26080
rect 50288 24992 50296 25056
rect 50360 24992 50376 25056
rect 50440 24992 50456 25056
rect 50520 24992 50536 25056
rect 50600 24992 50608 25056
rect 50288 23968 50608 24992
rect 50288 23904 50296 23968
rect 50360 23904 50376 23968
rect 50440 23904 50456 23968
rect 50520 23904 50536 23968
rect 50600 23904 50608 23968
rect 50288 22880 50608 23904
rect 50288 22816 50296 22880
rect 50360 22816 50376 22880
rect 50440 22816 50456 22880
rect 50520 22816 50536 22880
rect 50600 22816 50608 22880
rect 50288 21792 50608 22816
rect 50288 21728 50296 21792
rect 50360 21728 50376 21792
rect 50440 21728 50456 21792
rect 50520 21728 50536 21792
rect 50600 21728 50608 21792
rect 50288 20894 50608 21728
rect 50288 20704 50330 20894
rect 50566 20704 50608 20894
rect 50288 20640 50296 20704
rect 50360 20640 50376 20658
rect 50440 20640 50456 20658
rect 50520 20640 50536 20658
rect 50600 20640 50608 20704
rect 50288 19616 50608 20640
rect 50288 19552 50296 19616
rect 50360 19552 50376 19616
rect 50440 19552 50456 19616
rect 50520 19552 50536 19616
rect 50600 19552 50608 19616
rect 50288 18528 50608 19552
rect 50288 18464 50296 18528
rect 50360 18464 50376 18528
rect 50440 18464 50456 18528
rect 50520 18464 50536 18528
rect 50600 18464 50608 18528
rect 50288 17440 50608 18464
rect 50288 17376 50296 17440
rect 50360 17376 50376 17440
rect 50440 17376 50456 17440
rect 50520 17376 50536 17440
rect 50600 17376 50608 17440
rect 50288 16352 50608 17376
rect 50288 16288 50296 16352
rect 50360 16288 50376 16352
rect 50440 16288 50456 16352
rect 50520 16288 50536 16352
rect 50600 16288 50608 16352
rect 50288 15264 50608 16288
rect 50288 15200 50296 15264
rect 50360 15200 50376 15264
rect 50440 15200 50456 15264
rect 50520 15200 50536 15264
rect 50600 15200 50608 15264
rect 50288 14176 50608 15200
rect 50288 14112 50296 14176
rect 50360 14112 50376 14176
rect 50440 14112 50456 14176
rect 50520 14112 50536 14176
rect 50600 14112 50608 14176
rect 50288 13088 50608 14112
rect 50288 13024 50296 13088
rect 50360 13024 50376 13088
rect 50440 13024 50456 13088
rect 50520 13024 50536 13088
rect 50600 13024 50608 13088
rect 50288 12000 50608 13024
rect 50288 11936 50296 12000
rect 50360 11936 50376 12000
rect 50440 11936 50456 12000
rect 50520 11936 50536 12000
rect 50600 11936 50608 12000
rect 50288 10912 50608 11936
rect 50288 10848 50296 10912
rect 50360 10848 50376 10912
rect 50440 10848 50456 10912
rect 50520 10848 50536 10912
rect 50600 10848 50608 10912
rect 50288 9824 50608 10848
rect 50288 9760 50296 9824
rect 50360 9760 50376 9824
rect 50440 9760 50456 9824
rect 50520 9760 50536 9824
rect 50600 9760 50608 9824
rect 50288 8736 50608 9760
rect 50288 8672 50296 8736
rect 50360 8672 50376 8736
rect 50440 8672 50456 8736
rect 50520 8672 50536 8736
rect 50600 8672 50608 8736
rect 50288 7648 50608 8672
rect 50288 7584 50296 7648
rect 50360 7584 50376 7648
rect 50440 7584 50456 7648
rect 50520 7584 50536 7648
rect 50600 7584 50608 7648
rect 50288 6560 50608 7584
rect 50288 6496 50296 6560
rect 50360 6496 50376 6560
rect 50440 6496 50456 6560
rect 50520 6496 50536 6560
rect 50600 6496 50608 6560
rect 50288 5472 50608 6496
rect 50288 5408 50296 5472
rect 50360 5408 50376 5472
rect 50440 5408 50456 5472
rect 50520 5408 50536 5472
rect 50600 5408 50608 5472
rect 50288 4384 50608 5408
rect 50288 4320 50296 4384
rect 50360 4320 50376 4384
rect 50440 4320 50456 4384
rect 50520 4320 50536 4384
rect 50600 4320 50608 4384
rect 50288 3296 50608 4320
rect 50288 3232 50296 3296
rect 50360 3232 50376 3296
rect 50440 3232 50456 3296
rect 50520 3232 50536 3296
rect 50600 3232 50608 3296
rect 50288 2208 50608 3232
rect 50288 2144 50296 2208
rect 50360 2144 50376 2208
rect 50440 2144 50456 2208
rect 50520 2144 50536 2208
rect 50600 2144 50608 2208
rect 50288 2128 50608 2144
rect 65648 116992 65968 117552
rect 65648 116928 65656 116992
rect 65720 116928 65736 116992
rect 65800 116928 65816 116992
rect 65880 116928 65896 116992
rect 65960 116928 65968 116992
rect 65648 115904 65968 116928
rect 65648 115840 65656 115904
rect 65720 115840 65736 115904
rect 65800 115840 65816 115904
rect 65880 115840 65896 115904
rect 65960 115840 65968 115904
rect 65648 114816 65968 115840
rect 65648 114752 65656 114816
rect 65720 114752 65736 114816
rect 65800 114752 65816 114816
rect 65880 114752 65896 114816
rect 65960 114752 65968 114816
rect 65648 113728 65968 114752
rect 65648 113664 65656 113728
rect 65720 113664 65736 113728
rect 65800 113664 65816 113728
rect 65880 113664 65896 113728
rect 65960 113664 65968 113728
rect 65648 112640 65968 113664
rect 65648 112576 65656 112640
rect 65720 112576 65736 112640
rect 65800 112576 65816 112640
rect 65880 112576 65896 112640
rect 65960 112576 65968 112640
rect 65648 111552 65968 112576
rect 65648 111488 65656 111552
rect 65720 111488 65736 111552
rect 65800 111488 65816 111552
rect 65880 111488 65896 111552
rect 65960 111488 65968 111552
rect 65648 110464 65968 111488
rect 65648 110400 65656 110464
rect 65720 110400 65736 110464
rect 65800 110400 65816 110464
rect 65880 110400 65896 110464
rect 65960 110400 65968 110464
rect 65648 109376 65968 110400
rect 65648 109312 65656 109376
rect 65720 109312 65736 109376
rect 65800 109312 65816 109376
rect 65880 109312 65896 109376
rect 65960 109312 65968 109376
rect 65648 108288 65968 109312
rect 65648 108224 65656 108288
rect 65720 108224 65736 108288
rect 65800 108224 65816 108288
rect 65880 108224 65896 108288
rect 65960 108224 65968 108288
rect 65648 107200 65968 108224
rect 65648 107136 65656 107200
rect 65720 107136 65736 107200
rect 65800 107136 65816 107200
rect 65880 107136 65896 107200
rect 65960 107136 65968 107200
rect 65648 106112 65968 107136
rect 65648 106048 65656 106112
rect 65720 106048 65736 106112
rect 65800 106048 65816 106112
rect 65880 106048 65896 106112
rect 65960 106048 65968 106112
rect 65648 105024 65968 106048
rect 65648 104960 65656 105024
rect 65720 104960 65736 105024
rect 65800 104960 65816 105024
rect 65880 104960 65896 105024
rect 65960 104960 65968 105024
rect 65648 103936 65968 104960
rect 65648 103872 65656 103936
rect 65720 103872 65736 103936
rect 65800 103872 65816 103936
rect 65880 103872 65896 103936
rect 65960 103872 65968 103936
rect 65648 102848 65968 103872
rect 65648 102784 65656 102848
rect 65720 102784 65736 102848
rect 65800 102784 65816 102848
rect 65880 102784 65896 102848
rect 65960 102784 65968 102848
rect 65648 101760 65968 102784
rect 65648 101696 65656 101760
rect 65720 101696 65736 101760
rect 65800 101696 65816 101760
rect 65880 101696 65896 101760
rect 65960 101696 65968 101760
rect 65648 100672 65968 101696
rect 65648 100608 65656 100672
rect 65720 100608 65736 100672
rect 65800 100608 65816 100672
rect 65880 100608 65896 100672
rect 65960 100608 65968 100672
rect 65648 99584 65968 100608
rect 65648 99520 65656 99584
rect 65720 99520 65736 99584
rect 65800 99520 65816 99584
rect 65880 99520 65896 99584
rect 65960 99520 65968 99584
rect 65648 98496 65968 99520
rect 65648 98432 65656 98496
rect 65720 98432 65736 98496
rect 65800 98432 65816 98496
rect 65880 98432 65896 98496
rect 65960 98432 65968 98496
rect 65648 97484 65968 98432
rect 65648 97408 65690 97484
rect 65926 97408 65968 97484
rect 65648 97344 65656 97408
rect 65960 97344 65968 97408
rect 65648 97248 65690 97344
rect 65926 97248 65968 97344
rect 65648 96320 65968 97248
rect 65648 96256 65656 96320
rect 65720 96256 65736 96320
rect 65800 96256 65816 96320
rect 65880 96256 65896 96320
rect 65960 96256 65968 96320
rect 65648 95232 65968 96256
rect 65648 95168 65656 95232
rect 65720 95168 65736 95232
rect 65800 95168 65816 95232
rect 65880 95168 65896 95232
rect 65960 95168 65968 95232
rect 65648 94144 65968 95168
rect 65648 94080 65656 94144
rect 65720 94080 65736 94144
rect 65800 94080 65816 94144
rect 65880 94080 65896 94144
rect 65960 94080 65968 94144
rect 65648 93056 65968 94080
rect 65648 92992 65656 93056
rect 65720 92992 65736 93056
rect 65800 92992 65816 93056
rect 65880 92992 65896 93056
rect 65960 92992 65968 93056
rect 65648 91968 65968 92992
rect 65648 91904 65656 91968
rect 65720 91904 65736 91968
rect 65800 91904 65816 91968
rect 65880 91904 65896 91968
rect 65960 91904 65968 91968
rect 65648 90880 65968 91904
rect 65648 90816 65656 90880
rect 65720 90816 65736 90880
rect 65800 90816 65816 90880
rect 65880 90816 65896 90880
rect 65960 90816 65968 90880
rect 65648 89792 65968 90816
rect 65648 89728 65656 89792
rect 65720 89728 65736 89792
rect 65800 89728 65816 89792
rect 65880 89728 65896 89792
rect 65960 89728 65968 89792
rect 65648 88704 65968 89728
rect 65648 88640 65656 88704
rect 65720 88640 65736 88704
rect 65800 88640 65816 88704
rect 65880 88640 65896 88704
rect 65960 88640 65968 88704
rect 65648 87616 65968 88640
rect 65648 87552 65656 87616
rect 65720 87552 65736 87616
rect 65800 87552 65816 87616
rect 65880 87552 65896 87616
rect 65960 87552 65968 87616
rect 65648 86528 65968 87552
rect 65648 86464 65656 86528
rect 65720 86464 65736 86528
rect 65800 86464 65816 86528
rect 65880 86464 65896 86528
rect 65960 86464 65968 86528
rect 65648 85440 65968 86464
rect 65648 85376 65656 85440
rect 65720 85376 65736 85440
rect 65800 85376 65816 85440
rect 65880 85376 65896 85440
rect 65960 85376 65968 85440
rect 65648 84352 65968 85376
rect 65648 84288 65656 84352
rect 65720 84288 65736 84352
rect 65800 84288 65816 84352
rect 65880 84288 65896 84352
rect 65960 84288 65968 84352
rect 65648 83264 65968 84288
rect 65648 83200 65656 83264
rect 65720 83200 65736 83264
rect 65800 83200 65816 83264
rect 65880 83200 65896 83264
rect 65960 83200 65968 83264
rect 65648 82176 65968 83200
rect 65648 82112 65656 82176
rect 65720 82112 65736 82176
rect 65800 82112 65816 82176
rect 65880 82112 65896 82176
rect 65960 82112 65968 82176
rect 65648 81088 65968 82112
rect 65648 81024 65656 81088
rect 65720 81024 65736 81088
rect 65800 81024 65816 81088
rect 65880 81024 65896 81088
rect 65960 81024 65968 81088
rect 65648 80000 65968 81024
rect 65648 79936 65656 80000
rect 65720 79936 65736 80000
rect 65800 79936 65816 80000
rect 65880 79936 65896 80000
rect 65960 79936 65968 80000
rect 65648 78912 65968 79936
rect 65648 78848 65656 78912
rect 65720 78848 65736 78912
rect 65800 78848 65816 78912
rect 65880 78848 65896 78912
rect 65960 78848 65968 78912
rect 65648 77824 65968 78848
rect 65648 77760 65656 77824
rect 65720 77760 65736 77824
rect 65800 77760 65816 77824
rect 65880 77760 65896 77824
rect 65960 77760 65968 77824
rect 65648 76736 65968 77760
rect 65648 76672 65656 76736
rect 65720 76672 65736 76736
rect 65800 76672 65816 76736
rect 65880 76672 65896 76736
rect 65960 76672 65968 76736
rect 65648 75648 65968 76672
rect 65648 75584 65656 75648
rect 65720 75584 65736 75648
rect 65800 75584 65816 75648
rect 65880 75584 65896 75648
rect 65960 75584 65968 75648
rect 65648 74560 65968 75584
rect 65648 74496 65656 74560
rect 65720 74496 65736 74560
rect 65800 74496 65816 74560
rect 65880 74496 65896 74560
rect 65960 74496 65968 74560
rect 65648 73472 65968 74496
rect 65648 73408 65656 73472
rect 65720 73408 65736 73472
rect 65800 73408 65816 73472
rect 65880 73408 65896 73472
rect 65960 73408 65968 73472
rect 65648 72384 65968 73408
rect 65648 72320 65656 72384
rect 65720 72320 65736 72384
rect 65800 72320 65816 72384
rect 65880 72320 65896 72384
rect 65960 72320 65968 72384
rect 65648 71296 65968 72320
rect 65648 71232 65656 71296
rect 65720 71232 65736 71296
rect 65800 71232 65816 71296
rect 65880 71232 65896 71296
rect 65960 71232 65968 71296
rect 65648 70208 65968 71232
rect 65648 70144 65656 70208
rect 65720 70144 65736 70208
rect 65800 70144 65816 70208
rect 65880 70144 65896 70208
rect 65960 70144 65968 70208
rect 65648 69120 65968 70144
rect 65648 69056 65656 69120
rect 65720 69056 65736 69120
rect 65800 69056 65816 69120
rect 65880 69056 65896 69120
rect 65960 69056 65968 69120
rect 65648 68032 65968 69056
rect 65648 67968 65656 68032
rect 65720 67968 65736 68032
rect 65800 67968 65816 68032
rect 65880 67968 65896 68032
rect 65960 67968 65968 68032
rect 65648 66944 65968 67968
rect 65648 66880 65656 66944
rect 65720 66880 65736 66944
rect 65800 66880 65816 66944
rect 65880 66880 65896 66944
rect 65960 66880 65968 66944
rect 65648 66848 65968 66880
rect 65648 66612 65690 66848
rect 65926 66612 65968 66848
rect 65648 65856 65968 66612
rect 65648 65792 65656 65856
rect 65720 65792 65736 65856
rect 65800 65792 65816 65856
rect 65880 65792 65896 65856
rect 65960 65792 65968 65856
rect 65648 64768 65968 65792
rect 65648 64704 65656 64768
rect 65720 64704 65736 64768
rect 65800 64704 65816 64768
rect 65880 64704 65896 64768
rect 65960 64704 65968 64768
rect 65648 63680 65968 64704
rect 65648 63616 65656 63680
rect 65720 63616 65736 63680
rect 65800 63616 65816 63680
rect 65880 63616 65896 63680
rect 65960 63616 65968 63680
rect 65648 62592 65968 63616
rect 65648 62528 65656 62592
rect 65720 62528 65736 62592
rect 65800 62528 65816 62592
rect 65880 62528 65896 62592
rect 65960 62528 65968 62592
rect 65648 61504 65968 62528
rect 65648 61440 65656 61504
rect 65720 61440 65736 61504
rect 65800 61440 65816 61504
rect 65880 61440 65896 61504
rect 65960 61440 65968 61504
rect 65648 60416 65968 61440
rect 65648 60352 65656 60416
rect 65720 60352 65736 60416
rect 65800 60352 65816 60416
rect 65880 60352 65896 60416
rect 65960 60352 65968 60416
rect 65648 59328 65968 60352
rect 65648 59264 65656 59328
rect 65720 59264 65736 59328
rect 65800 59264 65816 59328
rect 65880 59264 65896 59328
rect 65960 59264 65968 59328
rect 65648 58240 65968 59264
rect 65648 58176 65656 58240
rect 65720 58176 65736 58240
rect 65800 58176 65816 58240
rect 65880 58176 65896 58240
rect 65960 58176 65968 58240
rect 65648 57152 65968 58176
rect 65648 57088 65656 57152
rect 65720 57088 65736 57152
rect 65800 57088 65816 57152
rect 65880 57088 65896 57152
rect 65960 57088 65968 57152
rect 65648 56064 65968 57088
rect 65648 56000 65656 56064
rect 65720 56000 65736 56064
rect 65800 56000 65816 56064
rect 65880 56000 65896 56064
rect 65960 56000 65968 56064
rect 65648 54976 65968 56000
rect 65648 54912 65656 54976
rect 65720 54912 65736 54976
rect 65800 54912 65816 54976
rect 65880 54912 65896 54976
rect 65960 54912 65968 54976
rect 65648 53888 65968 54912
rect 65648 53824 65656 53888
rect 65720 53824 65736 53888
rect 65800 53824 65816 53888
rect 65880 53824 65896 53888
rect 65960 53824 65968 53888
rect 65648 52800 65968 53824
rect 65648 52736 65656 52800
rect 65720 52736 65736 52800
rect 65800 52736 65816 52800
rect 65880 52736 65896 52800
rect 65960 52736 65968 52800
rect 65648 51712 65968 52736
rect 65648 51648 65656 51712
rect 65720 51648 65736 51712
rect 65800 51648 65816 51712
rect 65880 51648 65896 51712
rect 65960 51648 65968 51712
rect 65648 50624 65968 51648
rect 65648 50560 65656 50624
rect 65720 50560 65736 50624
rect 65800 50560 65816 50624
rect 65880 50560 65896 50624
rect 65960 50560 65968 50624
rect 65648 49536 65968 50560
rect 65648 49472 65656 49536
rect 65720 49472 65736 49536
rect 65800 49472 65816 49536
rect 65880 49472 65896 49536
rect 65960 49472 65968 49536
rect 65648 48448 65968 49472
rect 65648 48384 65656 48448
rect 65720 48384 65736 48448
rect 65800 48384 65816 48448
rect 65880 48384 65896 48448
rect 65960 48384 65968 48448
rect 65648 47360 65968 48384
rect 65648 47296 65656 47360
rect 65720 47296 65736 47360
rect 65800 47296 65816 47360
rect 65880 47296 65896 47360
rect 65960 47296 65968 47360
rect 65648 46272 65968 47296
rect 65648 46208 65656 46272
rect 65720 46208 65736 46272
rect 65800 46208 65816 46272
rect 65880 46208 65896 46272
rect 65960 46208 65968 46272
rect 65648 45184 65968 46208
rect 65648 45120 65656 45184
rect 65720 45120 65736 45184
rect 65800 45120 65816 45184
rect 65880 45120 65896 45184
rect 65960 45120 65968 45184
rect 65648 44096 65968 45120
rect 65648 44032 65656 44096
rect 65720 44032 65736 44096
rect 65800 44032 65816 44096
rect 65880 44032 65896 44096
rect 65960 44032 65968 44096
rect 65648 43008 65968 44032
rect 65648 42944 65656 43008
rect 65720 42944 65736 43008
rect 65800 42944 65816 43008
rect 65880 42944 65896 43008
rect 65960 42944 65968 43008
rect 65648 41920 65968 42944
rect 65648 41856 65656 41920
rect 65720 41856 65736 41920
rect 65800 41856 65816 41920
rect 65880 41856 65896 41920
rect 65960 41856 65968 41920
rect 65648 40832 65968 41856
rect 65648 40768 65656 40832
rect 65720 40768 65736 40832
rect 65800 40768 65816 40832
rect 65880 40768 65896 40832
rect 65960 40768 65968 40832
rect 65648 39744 65968 40768
rect 65648 39680 65656 39744
rect 65720 39680 65736 39744
rect 65800 39680 65816 39744
rect 65880 39680 65896 39744
rect 65960 39680 65968 39744
rect 65648 38656 65968 39680
rect 65648 38592 65656 38656
rect 65720 38592 65736 38656
rect 65800 38592 65816 38656
rect 65880 38592 65896 38656
rect 65960 38592 65968 38656
rect 65648 37568 65968 38592
rect 65648 37504 65656 37568
rect 65720 37504 65736 37568
rect 65800 37504 65816 37568
rect 65880 37504 65896 37568
rect 65960 37504 65968 37568
rect 65648 36480 65968 37504
rect 65648 36416 65656 36480
rect 65720 36416 65736 36480
rect 65800 36416 65816 36480
rect 65880 36416 65896 36480
rect 65960 36416 65968 36480
rect 65648 36212 65968 36416
rect 65648 35976 65690 36212
rect 65926 35976 65968 36212
rect 65648 35392 65968 35976
rect 65648 35328 65656 35392
rect 65720 35328 65736 35392
rect 65800 35328 65816 35392
rect 65880 35328 65896 35392
rect 65960 35328 65968 35392
rect 65648 34304 65968 35328
rect 65648 34240 65656 34304
rect 65720 34240 65736 34304
rect 65800 34240 65816 34304
rect 65880 34240 65896 34304
rect 65960 34240 65968 34304
rect 65648 33216 65968 34240
rect 65648 33152 65656 33216
rect 65720 33152 65736 33216
rect 65800 33152 65816 33216
rect 65880 33152 65896 33216
rect 65960 33152 65968 33216
rect 65648 32128 65968 33152
rect 65648 32064 65656 32128
rect 65720 32064 65736 32128
rect 65800 32064 65816 32128
rect 65880 32064 65896 32128
rect 65960 32064 65968 32128
rect 65648 31040 65968 32064
rect 65648 30976 65656 31040
rect 65720 30976 65736 31040
rect 65800 30976 65816 31040
rect 65880 30976 65896 31040
rect 65960 30976 65968 31040
rect 65648 29952 65968 30976
rect 65648 29888 65656 29952
rect 65720 29888 65736 29952
rect 65800 29888 65816 29952
rect 65880 29888 65896 29952
rect 65960 29888 65968 29952
rect 65648 28864 65968 29888
rect 65648 28800 65656 28864
rect 65720 28800 65736 28864
rect 65800 28800 65816 28864
rect 65880 28800 65896 28864
rect 65960 28800 65968 28864
rect 65648 27776 65968 28800
rect 65648 27712 65656 27776
rect 65720 27712 65736 27776
rect 65800 27712 65816 27776
rect 65880 27712 65896 27776
rect 65960 27712 65968 27776
rect 65648 26688 65968 27712
rect 65648 26624 65656 26688
rect 65720 26624 65736 26688
rect 65800 26624 65816 26688
rect 65880 26624 65896 26688
rect 65960 26624 65968 26688
rect 65648 25600 65968 26624
rect 65648 25536 65656 25600
rect 65720 25536 65736 25600
rect 65800 25536 65816 25600
rect 65880 25536 65896 25600
rect 65960 25536 65968 25600
rect 65648 24512 65968 25536
rect 65648 24448 65656 24512
rect 65720 24448 65736 24512
rect 65800 24448 65816 24512
rect 65880 24448 65896 24512
rect 65960 24448 65968 24512
rect 65648 23424 65968 24448
rect 65648 23360 65656 23424
rect 65720 23360 65736 23424
rect 65800 23360 65816 23424
rect 65880 23360 65896 23424
rect 65960 23360 65968 23424
rect 65648 22336 65968 23360
rect 65648 22272 65656 22336
rect 65720 22272 65736 22336
rect 65800 22272 65816 22336
rect 65880 22272 65896 22336
rect 65960 22272 65968 22336
rect 65648 21248 65968 22272
rect 65648 21184 65656 21248
rect 65720 21184 65736 21248
rect 65800 21184 65816 21248
rect 65880 21184 65896 21248
rect 65960 21184 65968 21248
rect 65648 20160 65968 21184
rect 65648 20096 65656 20160
rect 65720 20096 65736 20160
rect 65800 20096 65816 20160
rect 65880 20096 65896 20160
rect 65960 20096 65968 20160
rect 65648 19072 65968 20096
rect 65648 19008 65656 19072
rect 65720 19008 65736 19072
rect 65800 19008 65816 19072
rect 65880 19008 65896 19072
rect 65960 19008 65968 19072
rect 65648 17984 65968 19008
rect 65648 17920 65656 17984
rect 65720 17920 65736 17984
rect 65800 17920 65816 17984
rect 65880 17920 65896 17984
rect 65960 17920 65968 17984
rect 65648 16896 65968 17920
rect 65648 16832 65656 16896
rect 65720 16832 65736 16896
rect 65800 16832 65816 16896
rect 65880 16832 65896 16896
rect 65960 16832 65968 16896
rect 65648 15808 65968 16832
rect 65648 15744 65656 15808
rect 65720 15744 65736 15808
rect 65800 15744 65816 15808
rect 65880 15744 65896 15808
rect 65960 15744 65968 15808
rect 65648 14720 65968 15744
rect 65648 14656 65656 14720
rect 65720 14656 65736 14720
rect 65800 14656 65816 14720
rect 65880 14656 65896 14720
rect 65960 14656 65968 14720
rect 65648 13632 65968 14656
rect 65648 13568 65656 13632
rect 65720 13568 65736 13632
rect 65800 13568 65816 13632
rect 65880 13568 65896 13632
rect 65960 13568 65968 13632
rect 65648 12544 65968 13568
rect 65648 12480 65656 12544
rect 65720 12480 65736 12544
rect 65800 12480 65816 12544
rect 65880 12480 65896 12544
rect 65960 12480 65968 12544
rect 65648 11456 65968 12480
rect 65648 11392 65656 11456
rect 65720 11392 65736 11456
rect 65800 11392 65816 11456
rect 65880 11392 65896 11456
rect 65960 11392 65968 11456
rect 65648 10368 65968 11392
rect 65648 10304 65656 10368
rect 65720 10304 65736 10368
rect 65800 10304 65816 10368
rect 65880 10304 65896 10368
rect 65960 10304 65968 10368
rect 65648 9280 65968 10304
rect 65648 9216 65656 9280
rect 65720 9216 65736 9280
rect 65800 9216 65816 9280
rect 65880 9216 65896 9280
rect 65960 9216 65968 9280
rect 65648 8192 65968 9216
rect 65648 8128 65656 8192
rect 65720 8128 65736 8192
rect 65800 8128 65816 8192
rect 65880 8128 65896 8192
rect 65960 8128 65968 8192
rect 65648 7104 65968 8128
rect 65648 7040 65656 7104
rect 65720 7040 65736 7104
rect 65800 7040 65816 7104
rect 65880 7040 65896 7104
rect 65960 7040 65968 7104
rect 65648 6016 65968 7040
rect 65648 5952 65656 6016
rect 65720 5952 65736 6016
rect 65800 5952 65816 6016
rect 65880 5952 65896 6016
rect 65960 5952 65968 6016
rect 65648 5576 65968 5952
rect 65648 5340 65690 5576
rect 65926 5340 65968 5576
rect 65648 4928 65968 5340
rect 65648 4864 65656 4928
rect 65720 4864 65736 4928
rect 65800 4864 65816 4928
rect 65880 4864 65896 4928
rect 65960 4864 65968 4928
rect 65648 3840 65968 4864
rect 65648 3776 65656 3840
rect 65720 3776 65736 3840
rect 65800 3776 65816 3840
rect 65880 3776 65896 3840
rect 65960 3776 65968 3840
rect 65648 2752 65968 3776
rect 65648 2688 65656 2752
rect 65720 2688 65736 2752
rect 65800 2688 65816 2752
rect 65880 2688 65896 2752
rect 65960 2688 65968 2752
rect 65648 2128 65968 2688
<< via4 >>
rect 4250 97408 4486 97484
rect 4250 97344 4280 97408
rect 4280 97344 4296 97408
rect 4296 97344 4360 97408
rect 4360 97344 4376 97408
rect 4376 97344 4440 97408
rect 4440 97344 4456 97408
rect 4456 97344 4486 97408
rect 4250 97248 4486 97344
rect 4250 66612 4486 66848
rect 4250 35976 4486 36212
rect 4250 5340 4486 5576
rect 19610 112566 19846 112802
rect 19610 81930 19846 82166
rect 19610 51294 19846 51530
rect 19610 20704 19846 20894
rect 19610 20658 19640 20704
rect 19640 20658 19656 20704
rect 19656 20658 19720 20704
rect 19720 20658 19736 20704
rect 19736 20658 19800 20704
rect 19800 20658 19816 20704
rect 19816 20658 19846 20704
rect 34970 97408 35206 97484
rect 34970 97344 35000 97408
rect 35000 97344 35016 97408
rect 35016 97344 35080 97408
rect 35080 97344 35096 97408
rect 35096 97344 35160 97408
rect 35160 97344 35176 97408
rect 35176 97344 35206 97408
rect 34970 97248 35206 97344
rect 34970 66612 35206 66848
rect 34970 35976 35206 36212
rect 34970 5340 35206 5576
rect 50330 112566 50566 112802
rect 50330 81930 50566 82166
rect 50330 51294 50566 51530
rect 50330 20704 50566 20894
rect 50330 20658 50360 20704
rect 50360 20658 50376 20704
rect 50376 20658 50440 20704
rect 50440 20658 50456 20704
rect 50456 20658 50520 20704
rect 50520 20658 50536 20704
rect 50536 20658 50566 20704
rect 65690 97408 65926 97484
rect 65690 97344 65720 97408
rect 65720 97344 65736 97408
rect 65736 97344 65800 97408
rect 65800 97344 65816 97408
rect 65816 97344 65880 97408
rect 65880 97344 65896 97408
rect 65896 97344 65926 97408
rect 65690 97248 65926 97344
rect 65690 66612 65926 66848
rect 65690 35976 65926 36212
rect 65690 5340 65926 5576
<< metal5 >>
rect 1104 112802 78844 112844
rect 1104 112566 19610 112802
rect 19846 112566 50330 112802
rect 50566 112566 78844 112802
rect 1104 112524 78844 112566
rect 1104 97484 78844 97526
rect 1104 97248 4250 97484
rect 4486 97248 34970 97484
rect 35206 97248 65690 97484
rect 65926 97248 78844 97484
rect 1104 97206 78844 97248
rect 1104 82166 78844 82208
rect 1104 81930 19610 82166
rect 19846 81930 50330 82166
rect 50566 81930 78844 82166
rect 1104 81888 78844 81930
rect 1104 66848 78844 66890
rect 1104 66612 4250 66848
rect 4486 66612 34970 66848
rect 35206 66612 65690 66848
rect 65926 66612 78844 66848
rect 1104 66570 78844 66612
rect 1104 51530 78844 51572
rect 1104 51294 19610 51530
rect 19846 51294 50330 51530
rect 50566 51294 78844 51530
rect 1104 51252 78844 51294
rect 1104 36212 78844 36254
rect 1104 35976 4250 36212
rect 4486 35976 34970 36212
rect 35206 35976 65690 36212
rect 65926 35976 78844 36212
rect 1104 35934 78844 35976
rect 1104 20894 78844 20936
rect 1104 20658 19610 20894
rect 19846 20658 50330 20894
rect 50566 20658 78844 20894
rect 1104 20616 78844 20658
rect 1104 5576 78844 5618
rect 1104 5340 4250 5576
rect 4486 5340 34970 5576
rect 35206 5340 65690 5576
rect 65926 5340 78844 5576
rect 1104 5298 78844 5340
use sky130_fd_sc_hd__diode_2  ANTENNA_0 caravel_pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 2116 0 -1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1
timestamp 1644511149
transform 1 0 38548 0 -1 59840
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1644511149
transform 1 0 37720 0 1 59840
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1644511149
transform -1 0 39652 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp 1644511149
transform 1 0 35788 0 1 59840
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp 1644511149
transform 1 0 35236 0 -1 117504
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_6
timestamp 1644511149
transform -1 0 2116 0 1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_7
timestamp 1644511149
transform 1 0 66700 0 -1 117504
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_8
timestamp 1644511149
transform 1 0 77464 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_9
timestamp 1644511149
transform 1 0 2300 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_10
timestamp 1644511149
transform 1 0 74428 0 -1 117504
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_11
timestamp 1644511149
transform 1 0 77280 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_12
timestamp 1644511149
transform 1 0 73784 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_13
timestamp 1644511149
transform 1 0 77464 0 1 63104
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_14
timestamp 1644511149
transform -1 0 2116 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_15
timestamp 1644511149
transform 1 0 77280 0 -1 103360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_0_13 caravel_pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 2300 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25 caravel_pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3404 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_38
timestamp 1644511149
transform 1 0 4600 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50 caravel_pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 5704 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_57 caravel_pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 6348 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65 caravel_pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 7084 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_75
timestamp 1644511149
transform 1 0 8004 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_83
timestamp 1644511149
transform 1 0 8740 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_85
timestamp 1644511149
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_97
timestamp 1644511149
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_109
timestamp 1644511149
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_117
timestamp 1644511149
transform 1 0 11868 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_129
timestamp 1644511149
transform 1 0 12972 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_137
timestamp 1644511149
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_141
timestamp 1644511149
transform 1 0 14076 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_149
timestamp 1644511149
transform 1 0 14812 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_154
timestamp 1644511149
transform 1 0 15272 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_166 caravel_pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 16376 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_0_169
timestamp 1644511149
transform 1 0 16652 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_181 caravel_pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 17756 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_189
timestamp 1644511149
transform 1 0 18492 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_195
timestamp 1644511149
transform 1 0 19044 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_197
timestamp 1644511149
transform 1 0 19228 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_209
timestamp 1644511149
transform 1 0 20332 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_221
timestamp 1644511149
transform 1 0 21436 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_225
timestamp 1644511149
transform 1 0 21804 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_0_231
timestamp 1644511149
transform 1 0 22356 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_243
timestamp 1644511149
transform 1 0 23460 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_251
timestamp 1644511149
transform 1 0 24196 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_253
timestamp 1644511149
transform 1 0 24380 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_265
timestamp 1644511149
transform 1 0 25484 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_273
timestamp 1644511149
transform 1 0 26220 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_279
timestamp 1644511149
transform 1 0 26772 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_281
timestamp 1644511149
transform 1 0 26956 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_293
timestamp 1644511149
transform 1 0 28060 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_305
timestamp 1644511149
transform 1 0 29164 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_309
timestamp 1644511149
transform 1 0 29532 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_0_315
timestamp 1644511149
transform 1 0 30084 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_327
timestamp 1644511149
transform 1 0 31188 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_335
timestamp 1644511149
transform 1 0 31924 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_337
timestamp 1644511149
transform 1 0 32108 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_345
timestamp 1644511149
transform 1 0 32844 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_352
timestamp 1644511149
transform 1 0 33488 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_365
timestamp 1644511149
transform 1 0 34684 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_377
timestamp 1644511149
transform 1 0 35788 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_389
timestamp 1644511149
transform 1 0 36892 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_397
timestamp 1644511149
transform 1 0 37628 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_409
timestamp 1644511149
transform 1 0 38732 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_417
timestamp 1644511149
transform 1 0 39468 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_421
timestamp 1644511149
transform 1 0 39836 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_429
timestamp 1644511149
transform 1 0 40572 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_434
timestamp 1644511149
transform 1 0 41032 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_446
timestamp 1644511149
transform 1 0 42136 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_0_449
timestamp 1644511149
transform 1 0 42412 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_461
timestamp 1644511149
transform 1 0 43516 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_473
timestamp 1644511149
transform 1 0 44620 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_483
timestamp 1644511149
transform 1 0 45540 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_495
timestamp 1644511149
transform 1 0 46644 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_503
timestamp 1644511149
transform 1 0 47380 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_505
timestamp 1644511149
transform 1 0 47564 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_0_510
timestamp 1644511149
transform 1 0 48024 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_522
timestamp 1644511149
transform 1 0 49128 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_530
timestamp 1644511149
transform 1 0 49864 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_0_533
timestamp 1644511149
transform 1 0 50140 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_545
timestamp 1644511149
transform 1 0 51244 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_555
timestamp 1644511149
transform 1 0 52164 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_559
timestamp 1644511149
transform 1 0 52532 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_561
timestamp 1644511149
transform 1 0 52716 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_573
timestamp 1644511149
transform 1 0 53820 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_585
timestamp 1644511149
transform 1 0 54924 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_589
timestamp 1644511149
transform 1 0 55292 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_0_597
timestamp 1644511149
transform 1 0 56028 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_609
timestamp 1644511149
transform 1 0 57132 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_615
timestamp 1644511149
transform 1 0 57684 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_617
timestamp 1644511149
transform 1 0 57868 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_629
timestamp 1644511149
transform 1 0 58972 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_640
timestamp 1644511149
transform 1 0 59984 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_645
timestamp 1644511149
transform 1 0 60444 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_657
timestamp 1644511149
transform 1 0 61548 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_669
timestamp 1644511149
transform 1 0 62652 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_685
timestamp 1644511149
transform 1 0 64124 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_697
timestamp 1644511149
transform 1 0 65228 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_701
timestamp 1644511149
transform 1 0 65596 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_709
timestamp 1644511149
transform 1 0 66332 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_714
timestamp 1644511149
transform 1 0 66792 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_726
timestamp 1644511149
transform 1 0 67896 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_0_729
timestamp 1644511149
transform 1 0 68172 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_741
timestamp 1644511149
transform 1 0 69276 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_753
timestamp 1644511149
transform 1 0 70380 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_766
timestamp 1644511149
transform 1 0 71576 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_778
timestamp 1644511149
transform 1 0 72680 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_785
timestamp 1644511149
transform 1 0 73324 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_789
timestamp 1644511149
transform 1 0 73692 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_792
timestamp 1644511149
transform 1 0 73968 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_0_798
timestamp 1644511149
transform 1 0 74520 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_810
timestamp 1644511149
transform 1 0 75624 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_0_813
timestamp 1644511149
transform 1 0 75900 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_825
timestamp 1644511149
transform 1 0 77004 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_836
timestamp 1644511149
transform 1 0 78016 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_841
timestamp 1644511149
transform 1 0 78476 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_3
timestamp 1644511149
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_15
timestamp 1644511149
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_27
timestamp 1644511149
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_39
timestamp 1644511149
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_51
timestamp 1644511149
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1644511149
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_57
timestamp 1644511149
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_69
timestamp 1644511149
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_81
timestamp 1644511149
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_93
timestamp 1644511149
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_105
timestamp 1644511149
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 1644511149
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_113
timestamp 1644511149
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_125
timestamp 1644511149
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_137
timestamp 1644511149
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_149
timestamp 1644511149
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_161
timestamp 1644511149
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 1644511149
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_169
timestamp 1644511149
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_181
timestamp 1644511149
transform 1 0 17756 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_193
timestamp 1644511149
transform 1 0 18860 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_205
timestamp 1644511149
transform 1 0 19964 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_217
timestamp 1644511149
transform 1 0 21068 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_223
timestamp 1644511149
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_225
timestamp 1644511149
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_237
timestamp 1644511149
transform 1 0 22908 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_249
timestamp 1644511149
transform 1 0 24012 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_261
timestamp 1644511149
transform 1 0 25116 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_273
timestamp 1644511149
transform 1 0 26220 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_279
timestamp 1644511149
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_281
timestamp 1644511149
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_293
timestamp 1644511149
transform 1 0 28060 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_305
timestamp 1644511149
transform 1 0 29164 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_317
timestamp 1644511149
transform 1 0 30268 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_329
timestamp 1644511149
transform 1 0 31372 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_335
timestamp 1644511149
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_337
timestamp 1644511149
transform 1 0 32108 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_349
timestamp 1644511149
transform 1 0 33212 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_361
timestamp 1644511149
transform 1 0 34316 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_373
timestamp 1644511149
transform 1 0 35420 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_385
timestamp 1644511149
transform 1 0 36524 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_391
timestamp 1644511149
transform 1 0 37076 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_393
timestamp 1644511149
transform 1 0 37260 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_405
timestamp 1644511149
transform 1 0 38364 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_417
timestamp 1644511149
transform 1 0 39468 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_429
timestamp 1644511149
transform 1 0 40572 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_441
timestamp 1644511149
transform 1 0 41676 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_447
timestamp 1644511149
transform 1 0 42228 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_449
timestamp 1644511149
transform 1 0 42412 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_461
timestamp 1644511149
transform 1 0 43516 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_473
timestamp 1644511149
transform 1 0 44620 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_485
timestamp 1644511149
transform 1 0 45724 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_497
timestamp 1644511149
transform 1 0 46828 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_503
timestamp 1644511149
transform 1 0 47380 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_505
timestamp 1644511149
transform 1 0 47564 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_517
timestamp 1644511149
transform 1 0 48668 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_529
timestamp 1644511149
transform 1 0 49772 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_541
timestamp 1644511149
transform 1 0 50876 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_553
timestamp 1644511149
transform 1 0 51980 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_559
timestamp 1644511149
transform 1 0 52532 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_561
timestamp 1644511149
transform 1 0 52716 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_573
timestamp 1644511149
transform 1 0 53820 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_585
timestamp 1644511149
transform 1 0 54924 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_597
timestamp 1644511149
transform 1 0 56028 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_609
timestamp 1644511149
transform 1 0 57132 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_615
timestamp 1644511149
transform 1 0 57684 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_617
timestamp 1644511149
transform 1 0 57868 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_629
timestamp 1644511149
transform 1 0 58972 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_641
timestamp 1644511149
transform 1 0 60076 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_653
timestamp 1644511149
transform 1 0 61180 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_665
timestamp 1644511149
transform 1 0 62284 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_671
timestamp 1644511149
transform 1 0 62836 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_673
timestamp 1644511149
transform 1 0 63020 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_685
timestamp 1644511149
transform 1 0 64124 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_697
timestamp 1644511149
transform 1 0 65228 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_709
timestamp 1644511149
transform 1 0 66332 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_721
timestamp 1644511149
transform 1 0 67436 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_727
timestamp 1644511149
transform 1 0 67988 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_729
timestamp 1644511149
transform 1 0 68172 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_741
timestamp 1644511149
transform 1 0 69276 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_753
timestamp 1644511149
transform 1 0 70380 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_765
timestamp 1644511149
transform 1 0 71484 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_777
timestamp 1644511149
transform 1 0 72588 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_783
timestamp 1644511149
transform 1 0 73140 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_785
timestamp 1644511149
transform 1 0 73324 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_797
timestamp 1644511149
transform 1 0 74428 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_809
timestamp 1644511149
transform 1 0 75532 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_821
timestamp 1644511149
transform 1 0 76636 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_836
timestamp 1644511149
transform 1 0 78016 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_841
timestamp 1644511149
transform 1 0 78476 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_9
timestamp 1644511149
transform 1 0 1932 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_21
timestamp 1644511149
transform 1 0 3036 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1644511149
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_29
timestamp 1644511149
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_41
timestamp 1644511149
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_53
timestamp 1644511149
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_65
timestamp 1644511149
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp 1644511149
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1644511149
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_85
timestamp 1644511149
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_97
timestamp 1644511149
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_109
timestamp 1644511149
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_121
timestamp 1644511149
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_133
timestamp 1644511149
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 1644511149
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_141
timestamp 1644511149
transform 1 0 14076 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_149
timestamp 1644511149
transform 1 0 14812 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_153
timestamp 1644511149
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_165
timestamp 1644511149
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_177
timestamp 1644511149
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_189
timestamp 1644511149
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 1644511149
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_197
timestamp 1644511149
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_209
timestamp 1644511149
transform 1 0 20332 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_221
timestamp 1644511149
transform 1 0 21436 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_233
timestamp 1644511149
transform 1 0 22540 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_245
timestamp 1644511149
transform 1 0 23644 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_251
timestamp 1644511149
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_253
timestamp 1644511149
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_265
timestamp 1644511149
transform 1 0 25484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_277
timestamp 1644511149
transform 1 0 26588 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_289
timestamp 1644511149
transform 1 0 27692 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_301
timestamp 1644511149
transform 1 0 28796 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_307
timestamp 1644511149
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_309
timestamp 1644511149
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_321
timestamp 1644511149
transform 1 0 30636 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_333
timestamp 1644511149
transform 1 0 31740 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_345
timestamp 1644511149
transform 1 0 32844 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_357
timestamp 1644511149
transform 1 0 33948 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_363
timestamp 1644511149
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_365
timestamp 1644511149
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_377
timestamp 1644511149
transform 1 0 35788 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_389
timestamp 1644511149
transform 1 0 36892 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_401
timestamp 1644511149
transform 1 0 37996 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_413
timestamp 1644511149
transform 1 0 39100 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_419
timestamp 1644511149
transform 1 0 39652 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_421
timestamp 1644511149
transform 1 0 39836 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_429
timestamp 1644511149
transform 1 0 40572 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_437
timestamp 1644511149
transform 1 0 41308 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_444
timestamp 1644511149
transform 1 0 41952 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_456
timestamp 1644511149
transform 1 0 43056 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_468
timestamp 1644511149
transform 1 0 44160 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_2_477
timestamp 1644511149
transform 1 0 44988 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_489
timestamp 1644511149
transform 1 0 46092 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_501
timestamp 1644511149
transform 1 0 47196 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_513
timestamp 1644511149
transform 1 0 48300 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_525
timestamp 1644511149
transform 1 0 49404 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_531
timestamp 1644511149
transform 1 0 49956 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_533
timestamp 1644511149
transform 1 0 50140 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_545
timestamp 1644511149
transform 1 0 51244 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_557
timestamp 1644511149
transform 1 0 52348 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_569
timestamp 1644511149
transform 1 0 53452 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_581
timestamp 1644511149
transform 1 0 54556 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_587
timestamp 1644511149
transform 1 0 55108 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_589
timestamp 1644511149
transform 1 0 55292 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_601
timestamp 1644511149
transform 1 0 56396 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_613
timestamp 1644511149
transform 1 0 57500 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_625
timestamp 1644511149
transform 1 0 58604 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_637
timestamp 1644511149
transform 1 0 59708 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_643
timestamp 1644511149
transform 1 0 60260 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_645
timestamp 1644511149
transform 1 0 60444 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_657
timestamp 1644511149
transform 1 0 61548 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_669
timestamp 1644511149
transform 1 0 62652 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_681
timestamp 1644511149
transform 1 0 63756 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_693
timestamp 1644511149
transform 1 0 64860 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_699
timestamp 1644511149
transform 1 0 65412 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_701
timestamp 1644511149
transform 1 0 65596 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_713
timestamp 1644511149
transform 1 0 66700 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_725
timestamp 1644511149
transform 1 0 67804 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_737
timestamp 1644511149
transform 1 0 68908 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_749
timestamp 1644511149
transform 1 0 70012 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_755
timestamp 1644511149
transform 1 0 70564 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_757
timestamp 1644511149
transform 1 0 70748 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_769
timestamp 1644511149
transform 1 0 71852 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_781
timestamp 1644511149
transform 1 0 72956 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_793
timestamp 1644511149
transform 1 0 74060 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_805
timestamp 1644511149
transform 1 0 75164 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_811
timestamp 1644511149
transform 1 0 75716 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_813
timestamp 1644511149
transform 1 0 75900 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_825
timestamp 1644511149
transform 1 0 77004 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_837
timestamp 1644511149
transform 1 0 78108 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_841
timestamp 1644511149
transform 1 0 78476 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_3
timestamp 1644511149
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_15
timestamp 1644511149
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_27
timestamp 1644511149
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_39
timestamp 1644511149
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_51
timestamp 1644511149
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1644511149
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_57
timestamp 1644511149
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_69
timestamp 1644511149
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_81
timestamp 1644511149
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_93
timestamp 1644511149
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp 1644511149
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1644511149
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_113
timestamp 1644511149
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_125
timestamp 1644511149
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_137
timestamp 1644511149
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_149
timestamp 1644511149
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_161
timestamp 1644511149
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1644511149
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_169
timestamp 1644511149
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_181
timestamp 1644511149
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_193
timestamp 1644511149
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_205
timestamp 1644511149
transform 1 0 19964 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_217
timestamp 1644511149
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_223
timestamp 1644511149
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_225
timestamp 1644511149
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_237
timestamp 1644511149
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_249
timestamp 1644511149
transform 1 0 24012 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_261
timestamp 1644511149
transform 1 0 25116 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_273
timestamp 1644511149
transform 1 0 26220 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_279
timestamp 1644511149
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_281
timestamp 1644511149
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_293
timestamp 1644511149
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_305
timestamp 1644511149
transform 1 0 29164 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_317
timestamp 1644511149
transform 1 0 30268 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_329
timestamp 1644511149
transform 1 0 31372 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_335
timestamp 1644511149
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_337
timestamp 1644511149
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_349
timestamp 1644511149
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_361
timestamp 1644511149
transform 1 0 34316 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_373
timestamp 1644511149
transform 1 0 35420 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_385
timestamp 1644511149
transform 1 0 36524 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_391
timestamp 1644511149
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_393
timestamp 1644511149
transform 1 0 37260 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_405
timestamp 1644511149
transform 1 0 38364 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_417
timestamp 1644511149
transform 1 0 39468 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_429
timestamp 1644511149
transform 1 0 40572 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_441
timestamp 1644511149
transform 1 0 41676 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_447
timestamp 1644511149
transform 1 0 42228 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_449
timestamp 1644511149
transform 1 0 42412 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_461
timestamp 1644511149
transform 1 0 43516 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_473
timestamp 1644511149
transform 1 0 44620 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_485
timestamp 1644511149
transform 1 0 45724 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_497
timestamp 1644511149
transform 1 0 46828 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_503
timestamp 1644511149
transform 1 0 47380 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_505
timestamp 1644511149
transform 1 0 47564 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_517
timestamp 1644511149
transform 1 0 48668 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_529
timestamp 1644511149
transform 1 0 49772 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_541
timestamp 1644511149
transform 1 0 50876 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_553
timestamp 1644511149
transform 1 0 51980 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_559
timestamp 1644511149
transform 1 0 52532 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_561
timestamp 1644511149
transform 1 0 52716 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_573
timestamp 1644511149
transform 1 0 53820 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_585
timestamp 1644511149
transform 1 0 54924 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_597
timestamp 1644511149
transform 1 0 56028 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_609
timestamp 1644511149
transform 1 0 57132 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_615
timestamp 1644511149
transform 1 0 57684 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_617
timestamp 1644511149
transform 1 0 57868 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_629
timestamp 1644511149
transform 1 0 58972 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_641
timestamp 1644511149
transform 1 0 60076 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_653
timestamp 1644511149
transform 1 0 61180 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_665
timestamp 1644511149
transform 1 0 62284 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_671
timestamp 1644511149
transform 1 0 62836 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_673
timestamp 1644511149
transform 1 0 63020 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_685
timestamp 1644511149
transform 1 0 64124 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_697
timestamp 1644511149
transform 1 0 65228 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_709
timestamp 1644511149
transform 1 0 66332 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_721
timestamp 1644511149
transform 1 0 67436 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_727
timestamp 1644511149
transform 1 0 67988 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_729
timestamp 1644511149
transform 1 0 68172 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_741
timestamp 1644511149
transform 1 0 69276 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_753
timestamp 1644511149
transform 1 0 70380 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_765
timestamp 1644511149
transform 1 0 71484 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_777
timestamp 1644511149
transform 1 0 72588 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_783
timestamp 1644511149
transform 1 0 73140 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_785
timestamp 1644511149
transform 1 0 73324 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_797
timestamp 1644511149
transform 1 0 74428 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_809
timestamp 1644511149
transform 1 0 75532 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_821
timestamp 1644511149
transform 1 0 76636 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_833
timestamp 1644511149
transform 1 0 77740 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_839
timestamp 1644511149
transform 1 0 78292 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_841
timestamp 1644511149
transform 1 0 78476 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_3
timestamp 1644511149
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_15
timestamp 1644511149
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1644511149
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_29
timestamp 1644511149
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_41
timestamp 1644511149
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_53
timestamp 1644511149
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_65
timestamp 1644511149
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 1644511149
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1644511149
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_85
timestamp 1644511149
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_97
timestamp 1644511149
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_109
timestamp 1644511149
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_121
timestamp 1644511149
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp 1644511149
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1644511149
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_141
timestamp 1644511149
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_153
timestamp 1644511149
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_165
timestamp 1644511149
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_177
timestamp 1644511149
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_189
timestamp 1644511149
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 1644511149
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_197
timestamp 1644511149
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_209
timestamp 1644511149
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_221
timestamp 1644511149
transform 1 0 21436 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_233
timestamp 1644511149
transform 1 0 22540 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_245
timestamp 1644511149
transform 1 0 23644 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_251
timestamp 1644511149
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_253
timestamp 1644511149
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_265
timestamp 1644511149
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_277
timestamp 1644511149
transform 1 0 26588 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_289
timestamp 1644511149
transform 1 0 27692 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_301
timestamp 1644511149
transform 1 0 28796 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_307
timestamp 1644511149
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_309
timestamp 1644511149
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_321
timestamp 1644511149
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_333
timestamp 1644511149
transform 1 0 31740 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_345
timestamp 1644511149
transform 1 0 32844 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_357
timestamp 1644511149
transform 1 0 33948 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_363
timestamp 1644511149
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_365
timestamp 1644511149
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_377
timestamp 1644511149
transform 1 0 35788 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_389
timestamp 1644511149
transform 1 0 36892 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_401
timestamp 1644511149
transform 1 0 37996 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_413
timestamp 1644511149
transform 1 0 39100 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_419
timestamp 1644511149
transform 1 0 39652 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_421
timestamp 1644511149
transform 1 0 39836 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_433
timestamp 1644511149
transform 1 0 40940 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_445
timestamp 1644511149
transform 1 0 42044 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_457
timestamp 1644511149
transform 1 0 43148 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_469
timestamp 1644511149
transform 1 0 44252 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_475
timestamp 1644511149
transform 1 0 44804 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_477
timestamp 1644511149
transform 1 0 44988 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_489
timestamp 1644511149
transform 1 0 46092 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_501
timestamp 1644511149
transform 1 0 47196 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_513
timestamp 1644511149
transform 1 0 48300 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_525
timestamp 1644511149
transform 1 0 49404 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_531
timestamp 1644511149
transform 1 0 49956 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_533
timestamp 1644511149
transform 1 0 50140 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_545
timestamp 1644511149
transform 1 0 51244 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_557
timestamp 1644511149
transform 1 0 52348 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_569
timestamp 1644511149
transform 1 0 53452 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_581
timestamp 1644511149
transform 1 0 54556 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_587
timestamp 1644511149
transform 1 0 55108 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_589
timestamp 1644511149
transform 1 0 55292 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_601
timestamp 1644511149
transform 1 0 56396 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_613
timestamp 1644511149
transform 1 0 57500 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_625
timestamp 1644511149
transform 1 0 58604 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_637
timestamp 1644511149
transform 1 0 59708 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_643
timestamp 1644511149
transform 1 0 60260 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_645
timestamp 1644511149
transform 1 0 60444 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_657
timestamp 1644511149
transform 1 0 61548 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_669
timestamp 1644511149
transform 1 0 62652 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_681
timestamp 1644511149
transform 1 0 63756 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_693
timestamp 1644511149
transform 1 0 64860 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_699
timestamp 1644511149
transform 1 0 65412 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_701
timestamp 1644511149
transform 1 0 65596 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_713
timestamp 1644511149
transform 1 0 66700 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_725
timestamp 1644511149
transform 1 0 67804 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_737
timestamp 1644511149
transform 1 0 68908 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_749
timestamp 1644511149
transform 1 0 70012 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_755
timestamp 1644511149
transform 1 0 70564 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_757
timestamp 1644511149
transform 1 0 70748 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_769
timestamp 1644511149
transform 1 0 71852 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_781
timestamp 1644511149
transform 1 0 72956 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_793
timestamp 1644511149
transform 1 0 74060 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_805
timestamp 1644511149
transform 1 0 75164 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_811
timestamp 1644511149
transform 1 0 75716 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_813
timestamp 1644511149
transform 1 0 75900 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_825
timestamp 1644511149
transform 1 0 77004 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_833
timestamp 1644511149
transform 1 0 77740 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_837
timestamp 1644511149
transform 1 0 78108 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_841
timestamp 1644511149
transform 1 0 78476 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_3
timestamp 1644511149
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_15
timestamp 1644511149
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_27
timestamp 1644511149
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_39
timestamp 1644511149
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_51
timestamp 1644511149
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1644511149
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_57
timestamp 1644511149
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_69
timestamp 1644511149
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_81
timestamp 1644511149
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_93
timestamp 1644511149
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1644511149
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1644511149
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_113
timestamp 1644511149
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_125
timestamp 1644511149
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_137
timestamp 1644511149
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_149
timestamp 1644511149
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 1644511149
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1644511149
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_169
timestamp 1644511149
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_181
timestamp 1644511149
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_193
timestamp 1644511149
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_205
timestamp 1644511149
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_217
timestamp 1644511149
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_223
timestamp 1644511149
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_225
timestamp 1644511149
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_237
timestamp 1644511149
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_249
timestamp 1644511149
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_261
timestamp 1644511149
transform 1 0 25116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_273
timestamp 1644511149
transform 1 0 26220 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_279
timestamp 1644511149
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_281
timestamp 1644511149
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_293
timestamp 1644511149
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_305
timestamp 1644511149
transform 1 0 29164 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_317
timestamp 1644511149
transform 1 0 30268 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_329
timestamp 1644511149
transform 1 0 31372 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_335
timestamp 1644511149
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_337
timestamp 1644511149
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_349
timestamp 1644511149
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_361
timestamp 1644511149
transform 1 0 34316 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_373
timestamp 1644511149
transform 1 0 35420 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_385
timestamp 1644511149
transform 1 0 36524 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_391
timestamp 1644511149
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_393
timestamp 1644511149
transform 1 0 37260 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_405
timestamp 1644511149
transform 1 0 38364 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_417
timestamp 1644511149
transform 1 0 39468 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_429
timestamp 1644511149
transform 1 0 40572 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_441
timestamp 1644511149
transform 1 0 41676 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_447
timestamp 1644511149
transform 1 0 42228 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_449
timestamp 1644511149
transform 1 0 42412 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_461
timestamp 1644511149
transform 1 0 43516 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_473
timestamp 1644511149
transform 1 0 44620 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_485
timestamp 1644511149
transform 1 0 45724 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_497
timestamp 1644511149
transform 1 0 46828 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_503
timestamp 1644511149
transform 1 0 47380 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_505
timestamp 1644511149
transform 1 0 47564 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_517
timestamp 1644511149
transform 1 0 48668 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_529
timestamp 1644511149
transform 1 0 49772 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_541
timestamp 1644511149
transform 1 0 50876 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_553
timestamp 1644511149
transform 1 0 51980 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_559
timestamp 1644511149
transform 1 0 52532 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_561
timestamp 1644511149
transform 1 0 52716 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_573
timestamp 1644511149
transform 1 0 53820 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_585
timestamp 1644511149
transform 1 0 54924 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_597
timestamp 1644511149
transform 1 0 56028 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_609
timestamp 1644511149
transform 1 0 57132 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_615
timestamp 1644511149
transform 1 0 57684 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_617
timestamp 1644511149
transform 1 0 57868 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_629
timestamp 1644511149
transform 1 0 58972 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_641
timestamp 1644511149
transform 1 0 60076 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_653
timestamp 1644511149
transform 1 0 61180 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_665
timestamp 1644511149
transform 1 0 62284 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_671
timestamp 1644511149
transform 1 0 62836 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_673
timestamp 1644511149
transform 1 0 63020 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_685
timestamp 1644511149
transform 1 0 64124 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_697
timestamp 1644511149
transform 1 0 65228 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_709
timestamp 1644511149
transform 1 0 66332 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_721
timestamp 1644511149
transform 1 0 67436 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_727
timestamp 1644511149
transform 1 0 67988 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_729
timestamp 1644511149
transform 1 0 68172 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_741
timestamp 1644511149
transform 1 0 69276 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_753
timestamp 1644511149
transform 1 0 70380 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_765
timestamp 1644511149
transform 1 0 71484 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_777
timestamp 1644511149
transform 1 0 72588 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_783
timestamp 1644511149
transform 1 0 73140 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_785
timestamp 1644511149
transform 1 0 73324 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_797
timestamp 1644511149
transform 1 0 74428 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_809
timestamp 1644511149
transform 1 0 75532 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_821
timestamp 1644511149
transform 1 0 76636 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_829
timestamp 1644511149
transform 1 0 77372 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_836
timestamp 1644511149
transform 1 0 78016 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_841
timestamp 1644511149
transform 1 0 78476 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_3
timestamp 1644511149
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_15
timestamp 1644511149
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1644511149
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_29
timestamp 1644511149
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_41
timestamp 1644511149
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_53
timestamp 1644511149
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_65
timestamp 1644511149
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1644511149
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1644511149
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_85
timestamp 1644511149
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_97
timestamp 1644511149
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_109
timestamp 1644511149
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_121
timestamp 1644511149
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1644511149
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1644511149
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_141
timestamp 1644511149
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_153
timestamp 1644511149
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_165
timestamp 1644511149
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_177
timestamp 1644511149
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_189
timestamp 1644511149
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1644511149
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_197
timestamp 1644511149
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_209
timestamp 1644511149
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_221
timestamp 1644511149
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_233
timestamp 1644511149
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_245
timestamp 1644511149
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp 1644511149
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_253
timestamp 1644511149
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_265
timestamp 1644511149
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_277
timestamp 1644511149
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_289
timestamp 1644511149
transform 1 0 27692 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_301
timestamp 1644511149
transform 1 0 28796 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_307
timestamp 1644511149
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_309
timestamp 1644511149
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_321
timestamp 1644511149
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_333
timestamp 1644511149
transform 1 0 31740 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_345
timestamp 1644511149
transform 1 0 32844 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_357
timestamp 1644511149
transform 1 0 33948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_363
timestamp 1644511149
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_365
timestamp 1644511149
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_377
timestamp 1644511149
transform 1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_389
timestamp 1644511149
transform 1 0 36892 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_401
timestamp 1644511149
transform 1 0 37996 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_413
timestamp 1644511149
transform 1 0 39100 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_419
timestamp 1644511149
transform 1 0 39652 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_421
timestamp 1644511149
transform 1 0 39836 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_433
timestamp 1644511149
transform 1 0 40940 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_445
timestamp 1644511149
transform 1 0 42044 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_457
timestamp 1644511149
transform 1 0 43148 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_469
timestamp 1644511149
transform 1 0 44252 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_475
timestamp 1644511149
transform 1 0 44804 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_477
timestamp 1644511149
transform 1 0 44988 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_489
timestamp 1644511149
transform 1 0 46092 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_501
timestamp 1644511149
transform 1 0 47196 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_513
timestamp 1644511149
transform 1 0 48300 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_525
timestamp 1644511149
transform 1 0 49404 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_531
timestamp 1644511149
transform 1 0 49956 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_533
timestamp 1644511149
transform 1 0 50140 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_545
timestamp 1644511149
transform 1 0 51244 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_557
timestamp 1644511149
transform 1 0 52348 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_569
timestamp 1644511149
transform 1 0 53452 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_581
timestamp 1644511149
transform 1 0 54556 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_587
timestamp 1644511149
transform 1 0 55108 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_589
timestamp 1644511149
transform 1 0 55292 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_601
timestamp 1644511149
transform 1 0 56396 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_613
timestamp 1644511149
transform 1 0 57500 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_625
timestamp 1644511149
transform 1 0 58604 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_637
timestamp 1644511149
transform 1 0 59708 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_643
timestamp 1644511149
transform 1 0 60260 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_645
timestamp 1644511149
transform 1 0 60444 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_657
timestamp 1644511149
transform 1 0 61548 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_669
timestamp 1644511149
transform 1 0 62652 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_681
timestamp 1644511149
transform 1 0 63756 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_693
timestamp 1644511149
transform 1 0 64860 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_699
timestamp 1644511149
transform 1 0 65412 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_701
timestamp 1644511149
transform 1 0 65596 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_713
timestamp 1644511149
transform 1 0 66700 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_725
timestamp 1644511149
transform 1 0 67804 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_737
timestamp 1644511149
transform 1 0 68908 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_749
timestamp 1644511149
transform 1 0 70012 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_755
timestamp 1644511149
transform 1 0 70564 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_757
timestamp 1644511149
transform 1 0 70748 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_769
timestamp 1644511149
transform 1 0 71852 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_781
timestamp 1644511149
transform 1 0 72956 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_793
timestamp 1644511149
transform 1 0 74060 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_805
timestamp 1644511149
transform 1 0 75164 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_811
timestamp 1644511149
transform 1 0 75716 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_813
timestamp 1644511149
transform 1 0 75900 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_825
timestamp 1644511149
transform 1 0 77004 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_837
timestamp 1644511149
transform 1 0 78108 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_841
timestamp 1644511149
transform 1 0 78476 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_3
timestamp 1644511149
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_15
timestamp 1644511149
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_27
timestamp 1644511149
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_39
timestamp 1644511149
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp 1644511149
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1644511149
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_57
timestamp 1644511149
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_69
timestamp 1644511149
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_81
timestamp 1644511149
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_93
timestamp 1644511149
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1644511149
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1644511149
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_113
timestamp 1644511149
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_125
timestamp 1644511149
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_137
timestamp 1644511149
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_149
timestamp 1644511149
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp 1644511149
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1644511149
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_169
timestamp 1644511149
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_181
timestamp 1644511149
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_193
timestamp 1644511149
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_205
timestamp 1644511149
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_217
timestamp 1644511149
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp 1644511149
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_225
timestamp 1644511149
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_237
timestamp 1644511149
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_249
timestamp 1644511149
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_261
timestamp 1644511149
transform 1 0 25116 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_273
timestamp 1644511149
transform 1 0 26220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_279
timestamp 1644511149
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_281
timestamp 1644511149
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_293
timestamp 1644511149
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_305
timestamp 1644511149
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_317
timestamp 1644511149
transform 1 0 30268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_329
timestamp 1644511149
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_335
timestamp 1644511149
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_337
timestamp 1644511149
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_349
timestamp 1644511149
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_361
timestamp 1644511149
transform 1 0 34316 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_373
timestamp 1644511149
transform 1 0 35420 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_385
timestamp 1644511149
transform 1 0 36524 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_391
timestamp 1644511149
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_393
timestamp 1644511149
transform 1 0 37260 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_405
timestamp 1644511149
transform 1 0 38364 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_417
timestamp 1644511149
transform 1 0 39468 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_429
timestamp 1644511149
transform 1 0 40572 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_441
timestamp 1644511149
transform 1 0 41676 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_447
timestamp 1644511149
transform 1 0 42228 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_449
timestamp 1644511149
transform 1 0 42412 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_461
timestamp 1644511149
transform 1 0 43516 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_473
timestamp 1644511149
transform 1 0 44620 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_485
timestamp 1644511149
transform 1 0 45724 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_497
timestamp 1644511149
transform 1 0 46828 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_503
timestamp 1644511149
transform 1 0 47380 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_505
timestamp 1644511149
transform 1 0 47564 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_517
timestamp 1644511149
transform 1 0 48668 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_529
timestamp 1644511149
transform 1 0 49772 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_541
timestamp 1644511149
transform 1 0 50876 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_553
timestamp 1644511149
transform 1 0 51980 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_559
timestamp 1644511149
transform 1 0 52532 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_561
timestamp 1644511149
transform 1 0 52716 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_573
timestamp 1644511149
transform 1 0 53820 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_585
timestamp 1644511149
transform 1 0 54924 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_597
timestamp 1644511149
transform 1 0 56028 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_609
timestamp 1644511149
transform 1 0 57132 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_615
timestamp 1644511149
transform 1 0 57684 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_617
timestamp 1644511149
transform 1 0 57868 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_629
timestamp 1644511149
transform 1 0 58972 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_641
timestamp 1644511149
transform 1 0 60076 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_653
timestamp 1644511149
transform 1 0 61180 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_665
timestamp 1644511149
transform 1 0 62284 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_671
timestamp 1644511149
transform 1 0 62836 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_673
timestamp 1644511149
transform 1 0 63020 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_685
timestamp 1644511149
transform 1 0 64124 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_697
timestamp 1644511149
transform 1 0 65228 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_709
timestamp 1644511149
transform 1 0 66332 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_721
timestamp 1644511149
transform 1 0 67436 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_727
timestamp 1644511149
transform 1 0 67988 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_729
timestamp 1644511149
transform 1 0 68172 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_741
timestamp 1644511149
transform 1 0 69276 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_753
timestamp 1644511149
transform 1 0 70380 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_765
timestamp 1644511149
transform 1 0 71484 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_777
timestamp 1644511149
transform 1 0 72588 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_783
timestamp 1644511149
transform 1 0 73140 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_785
timestamp 1644511149
transform 1 0 73324 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_797
timestamp 1644511149
transform 1 0 74428 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_809
timestamp 1644511149
transform 1 0 75532 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_821
timestamp 1644511149
transform 1 0 76636 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_833
timestamp 1644511149
transform 1 0 77740 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_839
timestamp 1644511149
transform 1 0 78292 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_841
timestamp 1644511149
transform 1 0 78476 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_3
timestamp 1644511149
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_15
timestamp 1644511149
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1644511149
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_29
timestamp 1644511149
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_41
timestamp 1644511149
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_53
timestamp 1644511149
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_65
timestamp 1644511149
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1644511149
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1644511149
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_85
timestamp 1644511149
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_97
timestamp 1644511149
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_109
timestamp 1644511149
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_121
timestamp 1644511149
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp 1644511149
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1644511149
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_141
timestamp 1644511149
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_153
timestamp 1644511149
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_165
timestamp 1644511149
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_177
timestamp 1644511149
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_189
timestamp 1644511149
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1644511149
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_197
timestamp 1644511149
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_209
timestamp 1644511149
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_221
timestamp 1644511149
transform 1 0 21436 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_233
timestamp 1644511149
transform 1 0 22540 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_245
timestamp 1644511149
transform 1 0 23644 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_251
timestamp 1644511149
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_253
timestamp 1644511149
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_265
timestamp 1644511149
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_277
timestamp 1644511149
transform 1 0 26588 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_289
timestamp 1644511149
transform 1 0 27692 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_301
timestamp 1644511149
transform 1 0 28796 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_307
timestamp 1644511149
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_309
timestamp 1644511149
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_321
timestamp 1644511149
transform 1 0 30636 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_333
timestamp 1644511149
transform 1 0 31740 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_345
timestamp 1644511149
transform 1 0 32844 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_357
timestamp 1644511149
transform 1 0 33948 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_363
timestamp 1644511149
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_365
timestamp 1644511149
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_377
timestamp 1644511149
transform 1 0 35788 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_389
timestamp 1644511149
transform 1 0 36892 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_401
timestamp 1644511149
transform 1 0 37996 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_413
timestamp 1644511149
transform 1 0 39100 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_419
timestamp 1644511149
transform 1 0 39652 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_421
timestamp 1644511149
transform 1 0 39836 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_433
timestamp 1644511149
transform 1 0 40940 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_445
timestamp 1644511149
transform 1 0 42044 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_457
timestamp 1644511149
transform 1 0 43148 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_469
timestamp 1644511149
transform 1 0 44252 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_475
timestamp 1644511149
transform 1 0 44804 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_477
timestamp 1644511149
transform 1 0 44988 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_489
timestamp 1644511149
transform 1 0 46092 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_501
timestamp 1644511149
transform 1 0 47196 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_513
timestamp 1644511149
transform 1 0 48300 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_525
timestamp 1644511149
transform 1 0 49404 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_531
timestamp 1644511149
transform 1 0 49956 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_533
timestamp 1644511149
transform 1 0 50140 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_545
timestamp 1644511149
transform 1 0 51244 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_557
timestamp 1644511149
transform 1 0 52348 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_569
timestamp 1644511149
transform 1 0 53452 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_581
timestamp 1644511149
transform 1 0 54556 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_587
timestamp 1644511149
transform 1 0 55108 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_589
timestamp 1644511149
transform 1 0 55292 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_601
timestamp 1644511149
transform 1 0 56396 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_613
timestamp 1644511149
transform 1 0 57500 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_625
timestamp 1644511149
transform 1 0 58604 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_637
timestamp 1644511149
transform 1 0 59708 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_643
timestamp 1644511149
transform 1 0 60260 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_645
timestamp 1644511149
transform 1 0 60444 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_657
timestamp 1644511149
transform 1 0 61548 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_669
timestamp 1644511149
transform 1 0 62652 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_681
timestamp 1644511149
transform 1 0 63756 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_693
timestamp 1644511149
transform 1 0 64860 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_699
timestamp 1644511149
transform 1 0 65412 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_701
timestamp 1644511149
transform 1 0 65596 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_713
timestamp 1644511149
transform 1 0 66700 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_725
timestamp 1644511149
transform 1 0 67804 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_737
timestamp 1644511149
transform 1 0 68908 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_749
timestamp 1644511149
transform 1 0 70012 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_755
timestamp 1644511149
transform 1 0 70564 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_757
timestamp 1644511149
transform 1 0 70748 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_769
timestamp 1644511149
transform 1 0 71852 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_781
timestamp 1644511149
transform 1 0 72956 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_793
timestamp 1644511149
transform 1 0 74060 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_805
timestamp 1644511149
transform 1 0 75164 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_811
timestamp 1644511149
transform 1 0 75716 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_813
timestamp 1644511149
transform 1 0 75900 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_825
timestamp 1644511149
transform 1 0 77004 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_837
timestamp 1644511149
transform 1 0 78108 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_841
timestamp 1644511149
transform 1 0 78476 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_3
timestamp 1644511149
transform 1 0 1380 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_11
timestamp 1644511149
transform 1 0 2116 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_15
timestamp 1644511149
transform 1 0 2484 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_20
timestamp 1644511149
transform 1 0 2944 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_32
timestamp 1644511149
transform 1 0 4048 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_44
timestamp 1644511149
transform 1 0 5152 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_57
timestamp 1644511149
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_69
timestamp 1644511149
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_81
timestamp 1644511149
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_93
timestamp 1644511149
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp 1644511149
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1644511149
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_113
timestamp 1644511149
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_125
timestamp 1644511149
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_137
timestamp 1644511149
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_149
timestamp 1644511149
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_161
timestamp 1644511149
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1644511149
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_169
timestamp 1644511149
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_181
timestamp 1644511149
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_193
timestamp 1644511149
transform 1 0 18860 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_205
timestamp 1644511149
transform 1 0 19964 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_217
timestamp 1644511149
transform 1 0 21068 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_223
timestamp 1644511149
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_225
timestamp 1644511149
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_237
timestamp 1644511149
transform 1 0 22908 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_249
timestamp 1644511149
transform 1 0 24012 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_261
timestamp 1644511149
transform 1 0 25116 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_273
timestamp 1644511149
transform 1 0 26220 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_279
timestamp 1644511149
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_281
timestamp 1644511149
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_293
timestamp 1644511149
transform 1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_305
timestamp 1644511149
transform 1 0 29164 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_317
timestamp 1644511149
transform 1 0 30268 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_329
timestamp 1644511149
transform 1 0 31372 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_335
timestamp 1644511149
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_337
timestamp 1644511149
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_349
timestamp 1644511149
transform 1 0 33212 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_361
timestamp 1644511149
transform 1 0 34316 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_373
timestamp 1644511149
transform 1 0 35420 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_385
timestamp 1644511149
transform 1 0 36524 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_391
timestamp 1644511149
transform 1 0 37076 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_393
timestamp 1644511149
transform 1 0 37260 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_405
timestamp 1644511149
transform 1 0 38364 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_417
timestamp 1644511149
transform 1 0 39468 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_429
timestamp 1644511149
transform 1 0 40572 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_441
timestamp 1644511149
transform 1 0 41676 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_447
timestamp 1644511149
transform 1 0 42228 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_449
timestamp 1644511149
transform 1 0 42412 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_461
timestamp 1644511149
transform 1 0 43516 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_473
timestamp 1644511149
transform 1 0 44620 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_485
timestamp 1644511149
transform 1 0 45724 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_497
timestamp 1644511149
transform 1 0 46828 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_503
timestamp 1644511149
transform 1 0 47380 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_505
timestamp 1644511149
transform 1 0 47564 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_517
timestamp 1644511149
transform 1 0 48668 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_529
timestamp 1644511149
transform 1 0 49772 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_541
timestamp 1644511149
transform 1 0 50876 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_553
timestamp 1644511149
transform 1 0 51980 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_559
timestamp 1644511149
transform 1 0 52532 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_561
timestamp 1644511149
transform 1 0 52716 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_573
timestamp 1644511149
transform 1 0 53820 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_585
timestamp 1644511149
transform 1 0 54924 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_597
timestamp 1644511149
transform 1 0 56028 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_609
timestamp 1644511149
transform 1 0 57132 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_615
timestamp 1644511149
transform 1 0 57684 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_617
timestamp 1644511149
transform 1 0 57868 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_629
timestamp 1644511149
transform 1 0 58972 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_641
timestamp 1644511149
transform 1 0 60076 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_653
timestamp 1644511149
transform 1 0 61180 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_665
timestamp 1644511149
transform 1 0 62284 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_671
timestamp 1644511149
transform 1 0 62836 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_673
timestamp 1644511149
transform 1 0 63020 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_685
timestamp 1644511149
transform 1 0 64124 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_697
timestamp 1644511149
transform 1 0 65228 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_709
timestamp 1644511149
transform 1 0 66332 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_721
timestamp 1644511149
transform 1 0 67436 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_727
timestamp 1644511149
transform 1 0 67988 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_729
timestamp 1644511149
transform 1 0 68172 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_741
timestamp 1644511149
transform 1 0 69276 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_753
timestamp 1644511149
transform 1 0 70380 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_765
timestamp 1644511149
transform 1 0 71484 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_777
timestamp 1644511149
transform 1 0 72588 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_783
timestamp 1644511149
transform 1 0 73140 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_785
timestamp 1644511149
transform 1 0 73324 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_797
timestamp 1644511149
transform 1 0 74428 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_809
timestamp 1644511149
transform 1 0 75532 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_821
timestamp 1644511149
transform 1 0 76636 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_833
timestamp 1644511149
transform 1 0 77740 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_839
timestamp 1644511149
transform 1 0 78292 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_841
timestamp 1644511149
transform 1 0 78476 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_7
timestamp 1644511149
transform 1 0 1748 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_19
timestamp 1644511149
transform 1 0 2852 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1644511149
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_29
timestamp 1644511149
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_41
timestamp 1644511149
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_53
timestamp 1644511149
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_65
timestamp 1644511149
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 1644511149
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1644511149
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_85
timestamp 1644511149
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_97
timestamp 1644511149
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_109
timestamp 1644511149
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_121
timestamp 1644511149
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_133
timestamp 1644511149
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1644511149
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_141
timestamp 1644511149
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_153
timestamp 1644511149
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_165
timestamp 1644511149
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_177
timestamp 1644511149
transform 1 0 17388 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_189
timestamp 1644511149
transform 1 0 18492 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_195
timestamp 1644511149
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_197
timestamp 1644511149
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_209
timestamp 1644511149
transform 1 0 20332 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_221
timestamp 1644511149
transform 1 0 21436 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_233
timestamp 1644511149
transform 1 0 22540 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_245
timestamp 1644511149
transform 1 0 23644 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_251
timestamp 1644511149
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_253
timestamp 1644511149
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_265
timestamp 1644511149
transform 1 0 25484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_277
timestamp 1644511149
transform 1 0 26588 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_289
timestamp 1644511149
transform 1 0 27692 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_301
timestamp 1644511149
transform 1 0 28796 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_307
timestamp 1644511149
transform 1 0 29348 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_309
timestamp 1644511149
transform 1 0 29532 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_321
timestamp 1644511149
transform 1 0 30636 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_333
timestamp 1644511149
transform 1 0 31740 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_345
timestamp 1644511149
transform 1 0 32844 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_357
timestamp 1644511149
transform 1 0 33948 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_363
timestamp 1644511149
transform 1 0 34500 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_365
timestamp 1644511149
transform 1 0 34684 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_377
timestamp 1644511149
transform 1 0 35788 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_389
timestamp 1644511149
transform 1 0 36892 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_401
timestamp 1644511149
transform 1 0 37996 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_413
timestamp 1644511149
transform 1 0 39100 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_419
timestamp 1644511149
transform 1 0 39652 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_421
timestamp 1644511149
transform 1 0 39836 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_433
timestamp 1644511149
transform 1 0 40940 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_445
timestamp 1644511149
transform 1 0 42044 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_457
timestamp 1644511149
transform 1 0 43148 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_469
timestamp 1644511149
transform 1 0 44252 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_475
timestamp 1644511149
transform 1 0 44804 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_477
timestamp 1644511149
transform 1 0 44988 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_489
timestamp 1644511149
transform 1 0 46092 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_501
timestamp 1644511149
transform 1 0 47196 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_513
timestamp 1644511149
transform 1 0 48300 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_525
timestamp 1644511149
transform 1 0 49404 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_531
timestamp 1644511149
transform 1 0 49956 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_533
timestamp 1644511149
transform 1 0 50140 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_545
timestamp 1644511149
transform 1 0 51244 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_557
timestamp 1644511149
transform 1 0 52348 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_569
timestamp 1644511149
transform 1 0 53452 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_581
timestamp 1644511149
transform 1 0 54556 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_587
timestamp 1644511149
transform 1 0 55108 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_589
timestamp 1644511149
transform 1 0 55292 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_601
timestamp 1644511149
transform 1 0 56396 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_613
timestamp 1644511149
transform 1 0 57500 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_625
timestamp 1644511149
transform 1 0 58604 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_637
timestamp 1644511149
transform 1 0 59708 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_643
timestamp 1644511149
transform 1 0 60260 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_645
timestamp 1644511149
transform 1 0 60444 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_657
timestamp 1644511149
transform 1 0 61548 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_669
timestamp 1644511149
transform 1 0 62652 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_681
timestamp 1644511149
transform 1 0 63756 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_693
timestamp 1644511149
transform 1 0 64860 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_699
timestamp 1644511149
transform 1 0 65412 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_701
timestamp 1644511149
transform 1 0 65596 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_713
timestamp 1644511149
transform 1 0 66700 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_725
timestamp 1644511149
transform 1 0 67804 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_737
timestamp 1644511149
transform 1 0 68908 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_749
timestamp 1644511149
transform 1 0 70012 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_755
timestamp 1644511149
transform 1 0 70564 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_757
timestamp 1644511149
transform 1 0 70748 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_769
timestamp 1644511149
transform 1 0 71852 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_781
timestamp 1644511149
transform 1 0 72956 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_793
timestamp 1644511149
transform 1 0 74060 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_805
timestamp 1644511149
transform 1 0 75164 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_811
timestamp 1644511149
transform 1 0 75716 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_813
timestamp 1644511149
transform 1 0 75900 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_825
timestamp 1644511149
transform 1 0 77004 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_837
timestamp 1644511149
transform 1 0 78108 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_841
timestamp 1644511149
transform 1 0 78476 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_3
timestamp 1644511149
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_15
timestamp 1644511149
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_27
timestamp 1644511149
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_39
timestamp 1644511149
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_51
timestamp 1644511149
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1644511149
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_57
timestamp 1644511149
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_69
timestamp 1644511149
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_81
timestamp 1644511149
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_93
timestamp 1644511149
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_105
timestamp 1644511149
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1644511149
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_113
timestamp 1644511149
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_125
timestamp 1644511149
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_137
timestamp 1644511149
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_149
timestamp 1644511149
transform 1 0 14812 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_161
timestamp 1644511149
transform 1 0 15916 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp 1644511149
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_169
timestamp 1644511149
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_181
timestamp 1644511149
transform 1 0 17756 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_193
timestamp 1644511149
transform 1 0 18860 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_205
timestamp 1644511149
transform 1 0 19964 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_217
timestamp 1644511149
transform 1 0 21068 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_223
timestamp 1644511149
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_225
timestamp 1644511149
transform 1 0 21804 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_237
timestamp 1644511149
transform 1 0 22908 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_249
timestamp 1644511149
transform 1 0 24012 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_261
timestamp 1644511149
transform 1 0 25116 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_273
timestamp 1644511149
transform 1 0 26220 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_279
timestamp 1644511149
transform 1 0 26772 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_281
timestamp 1644511149
transform 1 0 26956 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_293
timestamp 1644511149
transform 1 0 28060 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_305
timestamp 1644511149
transform 1 0 29164 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_317
timestamp 1644511149
transform 1 0 30268 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_329
timestamp 1644511149
transform 1 0 31372 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_335
timestamp 1644511149
transform 1 0 31924 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_337
timestamp 1644511149
transform 1 0 32108 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_349
timestamp 1644511149
transform 1 0 33212 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_361
timestamp 1644511149
transform 1 0 34316 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_373
timestamp 1644511149
transform 1 0 35420 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_385
timestamp 1644511149
transform 1 0 36524 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_391
timestamp 1644511149
transform 1 0 37076 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_393
timestamp 1644511149
transform 1 0 37260 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_405
timestamp 1644511149
transform 1 0 38364 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_417
timestamp 1644511149
transform 1 0 39468 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_429
timestamp 1644511149
transform 1 0 40572 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_441
timestamp 1644511149
transform 1 0 41676 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_447
timestamp 1644511149
transform 1 0 42228 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_449
timestamp 1644511149
transform 1 0 42412 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_461
timestamp 1644511149
transform 1 0 43516 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_473
timestamp 1644511149
transform 1 0 44620 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_485
timestamp 1644511149
transform 1 0 45724 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_497
timestamp 1644511149
transform 1 0 46828 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_503
timestamp 1644511149
transform 1 0 47380 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_505
timestamp 1644511149
transform 1 0 47564 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_517
timestamp 1644511149
transform 1 0 48668 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_529
timestamp 1644511149
transform 1 0 49772 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_541
timestamp 1644511149
transform 1 0 50876 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_553
timestamp 1644511149
transform 1 0 51980 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_559
timestamp 1644511149
transform 1 0 52532 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_561
timestamp 1644511149
transform 1 0 52716 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_573
timestamp 1644511149
transform 1 0 53820 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_585
timestamp 1644511149
transform 1 0 54924 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_597
timestamp 1644511149
transform 1 0 56028 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_609
timestamp 1644511149
transform 1 0 57132 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_615
timestamp 1644511149
transform 1 0 57684 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_617
timestamp 1644511149
transform 1 0 57868 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_629
timestamp 1644511149
transform 1 0 58972 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_641
timestamp 1644511149
transform 1 0 60076 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_653
timestamp 1644511149
transform 1 0 61180 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_665
timestamp 1644511149
transform 1 0 62284 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_671
timestamp 1644511149
transform 1 0 62836 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_673
timestamp 1644511149
transform 1 0 63020 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_685
timestamp 1644511149
transform 1 0 64124 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_697
timestamp 1644511149
transform 1 0 65228 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_709
timestamp 1644511149
transform 1 0 66332 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_721
timestamp 1644511149
transform 1 0 67436 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_727
timestamp 1644511149
transform 1 0 67988 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_729
timestamp 1644511149
transform 1 0 68172 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_741
timestamp 1644511149
transform 1 0 69276 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_753
timestamp 1644511149
transform 1 0 70380 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_765
timestamp 1644511149
transform 1 0 71484 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_777
timestamp 1644511149
transform 1 0 72588 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_783
timestamp 1644511149
transform 1 0 73140 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_785
timestamp 1644511149
transform 1 0 73324 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_797
timestamp 1644511149
transform 1 0 74428 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_809
timestamp 1644511149
transform 1 0 75532 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_821
timestamp 1644511149
transform 1 0 76636 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_833
timestamp 1644511149
transform 1 0 77740 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_839
timestamp 1644511149
transform 1 0 78292 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_841
timestamp 1644511149
transform 1 0 78476 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_3
timestamp 1644511149
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_15
timestamp 1644511149
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1644511149
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_29
timestamp 1644511149
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_41
timestamp 1644511149
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_53
timestamp 1644511149
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_65
timestamp 1644511149
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1644511149
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1644511149
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_85
timestamp 1644511149
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_97
timestamp 1644511149
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_109
timestamp 1644511149
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_121
timestamp 1644511149
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_133
timestamp 1644511149
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1644511149
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_141
timestamp 1644511149
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_153
timestamp 1644511149
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_165
timestamp 1644511149
transform 1 0 16284 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_177
timestamp 1644511149
transform 1 0 17388 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_189
timestamp 1644511149
transform 1 0 18492 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_195
timestamp 1644511149
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_197
timestamp 1644511149
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_209
timestamp 1644511149
transform 1 0 20332 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_221
timestamp 1644511149
transform 1 0 21436 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_233
timestamp 1644511149
transform 1 0 22540 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_245
timestamp 1644511149
transform 1 0 23644 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_251
timestamp 1644511149
transform 1 0 24196 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_253
timestamp 1644511149
transform 1 0 24380 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_265
timestamp 1644511149
transform 1 0 25484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_277
timestamp 1644511149
transform 1 0 26588 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_289
timestamp 1644511149
transform 1 0 27692 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_301
timestamp 1644511149
transform 1 0 28796 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_307
timestamp 1644511149
transform 1 0 29348 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_309
timestamp 1644511149
transform 1 0 29532 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_321
timestamp 1644511149
transform 1 0 30636 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_333
timestamp 1644511149
transform 1 0 31740 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_345
timestamp 1644511149
transform 1 0 32844 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_357
timestamp 1644511149
transform 1 0 33948 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_363
timestamp 1644511149
transform 1 0 34500 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_365
timestamp 1644511149
transform 1 0 34684 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_377
timestamp 1644511149
transform 1 0 35788 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_389
timestamp 1644511149
transform 1 0 36892 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_401
timestamp 1644511149
transform 1 0 37996 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_413
timestamp 1644511149
transform 1 0 39100 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_419
timestamp 1644511149
transform 1 0 39652 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_421
timestamp 1644511149
transform 1 0 39836 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_433
timestamp 1644511149
transform 1 0 40940 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_445
timestamp 1644511149
transform 1 0 42044 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_457
timestamp 1644511149
transform 1 0 43148 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_469
timestamp 1644511149
transform 1 0 44252 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_475
timestamp 1644511149
transform 1 0 44804 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_477
timestamp 1644511149
transform 1 0 44988 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_489
timestamp 1644511149
transform 1 0 46092 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_501
timestamp 1644511149
transform 1 0 47196 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_513
timestamp 1644511149
transform 1 0 48300 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_525
timestamp 1644511149
transform 1 0 49404 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_531
timestamp 1644511149
transform 1 0 49956 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_533
timestamp 1644511149
transform 1 0 50140 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_545
timestamp 1644511149
transform 1 0 51244 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_557
timestamp 1644511149
transform 1 0 52348 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_569
timestamp 1644511149
transform 1 0 53452 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_581
timestamp 1644511149
transform 1 0 54556 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_587
timestamp 1644511149
transform 1 0 55108 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_589
timestamp 1644511149
transform 1 0 55292 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_601
timestamp 1644511149
transform 1 0 56396 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_613
timestamp 1644511149
transform 1 0 57500 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_625
timestamp 1644511149
transform 1 0 58604 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_637
timestamp 1644511149
transform 1 0 59708 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_643
timestamp 1644511149
transform 1 0 60260 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_645
timestamp 1644511149
transform 1 0 60444 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_657
timestamp 1644511149
transform 1 0 61548 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_669
timestamp 1644511149
transform 1 0 62652 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_681
timestamp 1644511149
transform 1 0 63756 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_693
timestamp 1644511149
transform 1 0 64860 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_699
timestamp 1644511149
transform 1 0 65412 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_701
timestamp 1644511149
transform 1 0 65596 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_713
timestamp 1644511149
transform 1 0 66700 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_725
timestamp 1644511149
transform 1 0 67804 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_737
timestamp 1644511149
transform 1 0 68908 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_749
timestamp 1644511149
transform 1 0 70012 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_755
timestamp 1644511149
transform 1 0 70564 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_757
timestamp 1644511149
transform 1 0 70748 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_769
timestamp 1644511149
transform 1 0 71852 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_781
timestamp 1644511149
transform 1 0 72956 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_793
timestamp 1644511149
transform 1 0 74060 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_805
timestamp 1644511149
transform 1 0 75164 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_811
timestamp 1644511149
transform 1 0 75716 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_813
timestamp 1644511149
transform 1 0 75900 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_825
timestamp 1644511149
transform 1 0 77004 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_829
timestamp 1644511149
transform 1 0 77372 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_832
timestamp 1644511149
transform 1 0 77648 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_838
timestamp 1644511149
transform 1 0 78200 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_3
timestamp 1644511149
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_15
timestamp 1644511149
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_27
timestamp 1644511149
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_39
timestamp 1644511149
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_51
timestamp 1644511149
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1644511149
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_57
timestamp 1644511149
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_69
timestamp 1644511149
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_81
timestamp 1644511149
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_93
timestamp 1644511149
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_105
timestamp 1644511149
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1644511149
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_113
timestamp 1644511149
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_125
timestamp 1644511149
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_137
timestamp 1644511149
transform 1 0 13708 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_149
timestamp 1644511149
transform 1 0 14812 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_161
timestamp 1644511149
transform 1 0 15916 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1644511149
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_169
timestamp 1644511149
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_181
timestamp 1644511149
transform 1 0 17756 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_193
timestamp 1644511149
transform 1 0 18860 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_205
timestamp 1644511149
transform 1 0 19964 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_217
timestamp 1644511149
transform 1 0 21068 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_223
timestamp 1644511149
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_225
timestamp 1644511149
transform 1 0 21804 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_237
timestamp 1644511149
transform 1 0 22908 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_249
timestamp 1644511149
transform 1 0 24012 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_261
timestamp 1644511149
transform 1 0 25116 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_273
timestamp 1644511149
transform 1 0 26220 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_279
timestamp 1644511149
transform 1 0 26772 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_281
timestamp 1644511149
transform 1 0 26956 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_293
timestamp 1644511149
transform 1 0 28060 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_305
timestamp 1644511149
transform 1 0 29164 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_317
timestamp 1644511149
transform 1 0 30268 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_329
timestamp 1644511149
transform 1 0 31372 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_335
timestamp 1644511149
transform 1 0 31924 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_337
timestamp 1644511149
transform 1 0 32108 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_349
timestamp 1644511149
transform 1 0 33212 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_361
timestamp 1644511149
transform 1 0 34316 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_373
timestamp 1644511149
transform 1 0 35420 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_385
timestamp 1644511149
transform 1 0 36524 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_391
timestamp 1644511149
transform 1 0 37076 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_393
timestamp 1644511149
transform 1 0 37260 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_405
timestamp 1644511149
transform 1 0 38364 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_417
timestamp 1644511149
transform 1 0 39468 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_429
timestamp 1644511149
transform 1 0 40572 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_441
timestamp 1644511149
transform 1 0 41676 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_447
timestamp 1644511149
transform 1 0 42228 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_449
timestamp 1644511149
transform 1 0 42412 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_461
timestamp 1644511149
transform 1 0 43516 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_473
timestamp 1644511149
transform 1 0 44620 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_485
timestamp 1644511149
transform 1 0 45724 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_497
timestamp 1644511149
transform 1 0 46828 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_503
timestamp 1644511149
transform 1 0 47380 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_505
timestamp 1644511149
transform 1 0 47564 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_517
timestamp 1644511149
transform 1 0 48668 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_529
timestamp 1644511149
transform 1 0 49772 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_541
timestamp 1644511149
transform 1 0 50876 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_553
timestamp 1644511149
transform 1 0 51980 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_559
timestamp 1644511149
transform 1 0 52532 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_561
timestamp 1644511149
transform 1 0 52716 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_573
timestamp 1644511149
transform 1 0 53820 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_585
timestamp 1644511149
transform 1 0 54924 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_597
timestamp 1644511149
transform 1 0 56028 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_609
timestamp 1644511149
transform 1 0 57132 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_615
timestamp 1644511149
transform 1 0 57684 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_617
timestamp 1644511149
transform 1 0 57868 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_629
timestamp 1644511149
transform 1 0 58972 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_641
timestamp 1644511149
transform 1 0 60076 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_653
timestamp 1644511149
transform 1 0 61180 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_665
timestamp 1644511149
transform 1 0 62284 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_671
timestamp 1644511149
transform 1 0 62836 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_673
timestamp 1644511149
transform 1 0 63020 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_685
timestamp 1644511149
transform 1 0 64124 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_697
timestamp 1644511149
transform 1 0 65228 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_709
timestamp 1644511149
transform 1 0 66332 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_721
timestamp 1644511149
transform 1 0 67436 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_727
timestamp 1644511149
transform 1 0 67988 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_729
timestamp 1644511149
transform 1 0 68172 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_741
timestamp 1644511149
transform 1 0 69276 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_753
timestamp 1644511149
transform 1 0 70380 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_765
timestamp 1644511149
transform 1 0 71484 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_777
timestamp 1644511149
transform 1 0 72588 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_783
timestamp 1644511149
transform 1 0 73140 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_785
timestamp 1644511149
transform 1 0 73324 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_797
timestamp 1644511149
transform 1 0 74428 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_809
timestamp 1644511149
transform 1 0 75532 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_821
timestamp 1644511149
transform 1 0 76636 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_833
timestamp 1644511149
transform 1 0 77740 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_839
timestamp 1644511149
transform 1 0 78292 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_841
timestamp 1644511149
transform 1 0 78476 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_3
timestamp 1644511149
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_15
timestamp 1644511149
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1644511149
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_29
timestamp 1644511149
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_41
timestamp 1644511149
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_53
timestamp 1644511149
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_65
timestamp 1644511149
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 1644511149
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1644511149
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_85
timestamp 1644511149
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_97
timestamp 1644511149
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_109
timestamp 1644511149
transform 1 0 11132 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_121
timestamp 1644511149
transform 1 0 12236 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_133
timestamp 1644511149
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1644511149
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_141
timestamp 1644511149
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_153
timestamp 1644511149
transform 1 0 15180 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_165
timestamp 1644511149
transform 1 0 16284 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_177
timestamp 1644511149
transform 1 0 17388 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_189
timestamp 1644511149
transform 1 0 18492 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_195
timestamp 1644511149
transform 1 0 19044 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_197
timestamp 1644511149
transform 1 0 19228 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_209
timestamp 1644511149
transform 1 0 20332 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_221
timestamp 1644511149
transform 1 0 21436 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_233
timestamp 1644511149
transform 1 0 22540 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_245
timestamp 1644511149
transform 1 0 23644 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_251
timestamp 1644511149
transform 1 0 24196 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_253
timestamp 1644511149
transform 1 0 24380 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_265
timestamp 1644511149
transform 1 0 25484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_277
timestamp 1644511149
transform 1 0 26588 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_289
timestamp 1644511149
transform 1 0 27692 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_301
timestamp 1644511149
transform 1 0 28796 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_307
timestamp 1644511149
transform 1 0 29348 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_309
timestamp 1644511149
transform 1 0 29532 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_321
timestamp 1644511149
transform 1 0 30636 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_333
timestamp 1644511149
transform 1 0 31740 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_345
timestamp 1644511149
transform 1 0 32844 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_357
timestamp 1644511149
transform 1 0 33948 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_363
timestamp 1644511149
transform 1 0 34500 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_365
timestamp 1644511149
transform 1 0 34684 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_377
timestamp 1644511149
transform 1 0 35788 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_389
timestamp 1644511149
transform 1 0 36892 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_401
timestamp 1644511149
transform 1 0 37996 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_413
timestamp 1644511149
transform 1 0 39100 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_419
timestamp 1644511149
transform 1 0 39652 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_421
timestamp 1644511149
transform 1 0 39836 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_433
timestamp 1644511149
transform 1 0 40940 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_445
timestamp 1644511149
transform 1 0 42044 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_457
timestamp 1644511149
transform 1 0 43148 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_469
timestamp 1644511149
transform 1 0 44252 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_475
timestamp 1644511149
transform 1 0 44804 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_477
timestamp 1644511149
transform 1 0 44988 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_489
timestamp 1644511149
transform 1 0 46092 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_501
timestamp 1644511149
transform 1 0 47196 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_513
timestamp 1644511149
transform 1 0 48300 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_525
timestamp 1644511149
transform 1 0 49404 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_531
timestamp 1644511149
transform 1 0 49956 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_533
timestamp 1644511149
transform 1 0 50140 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_545
timestamp 1644511149
transform 1 0 51244 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_557
timestamp 1644511149
transform 1 0 52348 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_569
timestamp 1644511149
transform 1 0 53452 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_581
timestamp 1644511149
transform 1 0 54556 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_587
timestamp 1644511149
transform 1 0 55108 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_589
timestamp 1644511149
transform 1 0 55292 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_601
timestamp 1644511149
transform 1 0 56396 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_613
timestamp 1644511149
transform 1 0 57500 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_625
timestamp 1644511149
transform 1 0 58604 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_637
timestamp 1644511149
transform 1 0 59708 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_643
timestamp 1644511149
transform 1 0 60260 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_645
timestamp 1644511149
transform 1 0 60444 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_657
timestamp 1644511149
transform 1 0 61548 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_669
timestamp 1644511149
transform 1 0 62652 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_681
timestamp 1644511149
transform 1 0 63756 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_693
timestamp 1644511149
transform 1 0 64860 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_699
timestamp 1644511149
transform 1 0 65412 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_701
timestamp 1644511149
transform 1 0 65596 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_713
timestamp 1644511149
transform 1 0 66700 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_725
timestamp 1644511149
transform 1 0 67804 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_737
timestamp 1644511149
transform 1 0 68908 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_749
timestamp 1644511149
transform 1 0 70012 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_755
timestamp 1644511149
transform 1 0 70564 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_757
timestamp 1644511149
transform 1 0 70748 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_769
timestamp 1644511149
transform 1 0 71852 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_781
timestamp 1644511149
transform 1 0 72956 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_793
timestamp 1644511149
transform 1 0 74060 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_805
timestamp 1644511149
transform 1 0 75164 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_811
timestamp 1644511149
transform 1 0 75716 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_813
timestamp 1644511149
transform 1 0 75900 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_825
timestamp 1644511149
transform 1 0 77004 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_838
timestamp 1644511149
transform 1 0 78200 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_15_3
timestamp 1644511149
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_15
timestamp 1644511149
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_27
timestamp 1644511149
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_39
timestamp 1644511149
transform 1 0 4692 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_51
timestamp 1644511149
transform 1 0 5796 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1644511149
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_57
timestamp 1644511149
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_69
timestamp 1644511149
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_81
timestamp 1644511149
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_93
timestamp 1644511149
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_105
timestamp 1644511149
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1644511149
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_113
timestamp 1644511149
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_125
timestamp 1644511149
transform 1 0 12604 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_137
timestamp 1644511149
transform 1 0 13708 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_149
timestamp 1644511149
transform 1 0 14812 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_161
timestamp 1644511149
transform 1 0 15916 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_167
timestamp 1644511149
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_169
timestamp 1644511149
transform 1 0 16652 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_181
timestamp 1644511149
transform 1 0 17756 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_193
timestamp 1644511149
transform 1 0 18860 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_205
timestamp 1644511149
transform 1 0 19964 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_217
timestamp 1644511149
transform 1 0 21068 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_223
timestamp 1644511149
transform 1 0 21620 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_225
timestamp 1644511149
transform 1 0 21804 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_237
timestamp 1644511149
transform 1 0 22908 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_249
timestamp 1644511149
transform 1 0 24012 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_261
timestamp 1644511149
transform 1 0 25116 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_273
timestamp 1644511149
transform 1 0 26220 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_279
timestamp 1644511149
transform 1 0 26772 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_281
timestamp 1644511149
transform 1 0 26956 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_293
timestamp 1644511149
transform 1 0 28060 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_305
timestamp 1644511149
transform 1 0 29164 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_317
timestamp 1644511149
transform 1 0 30268 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_329
timestamp 1644511149
transform 1 0 31372 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_335
timestamp 1644511149
transform 1 0 31924 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_337
timestamp 1644511149
transform 1 0 32108 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_349
timestamp 1644511149
transform 1 0 33212 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_361
timestamp 1644511149
transform 1 0 34316 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_373
timestamp 1644511149
transform 1 0 35420 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_385
timestamp 1644511149
transform 1 0 36524 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_391
timestamp 1644511149
transform 1 0 37076 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_393
timestamp 1644511149
transform 1 0 37260 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_405
timestamp 1644511149
transform 1 0 38364 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_417
timestamp 1644511149
transform 1 0 39468 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_429
timestamp 1644511149
transform 1 0 40572 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_441
timestamp 1644511149
transform 1 0 41676 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_447
timestamp 1644511149
transform 1 0 42228 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_449
timestamp 1644511149
transform 1 0 42412 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_461
timestamp 1644511149
transform 1 0 43516 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_473
timestamp 1644511149
transform 1 0 44620 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_485
timestamp 1644511149
transform 1 0 45724 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_497
timestamp 1644511149
transform 1 0 46828 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_503
timestamp 1644511149
transform 1 0 47380 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_505
timestamp 1644511149
transform 1 0 47564 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_517
timestamp 1644511149
transform 1 0 48668 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_529
timestamp 1644511149
transform 1 0 49772 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_541
timestamp 1644511149
transform 1 0 50876 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_553
timestamp 1644511149
transform 1 0 51980 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_559
timestamp 1644511149
transform 1 0 52532 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_561
timestamp 1644511149
transform 1 0 52716 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_573
timestamp 1644511149
transform 1 0 53820 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_585
timestamp 1644511149
transform 1 0 54924 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_597
timestamp 1644511149
transform 1 0 56028 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_609
timestamp 1644511149
transform 1 0 57132 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_615
timestamp 1644511149
transform 1 0 57684 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_617
timestamp 1644511149
transform 1 0 57868 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_629
timestamp 1644511149
transform 1 0 58972 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_641
timestamp 1644511149
transform 1 0 60076 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_653
timestamp 1644511149
transform 1 0 61180 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_665
timestamp 1644511149
transform 1 0 62284 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_671
timestamp 1644511149
transform 1 0 62836 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_673
timestamp 1644511149
transform 1 0 63020 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_685
timestamp 1644511149
transform 1 0 64124 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_697
timestamp 1644511149
transform 1 0 65228 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_709
timestamp 1644511149
transform 1 0 66332 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_721
timestamp 1644511149
transform 1 0 67436 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_727
timestamp 1644511149
transform 1 0 67988 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_729
timestamp 1644511149
transform 1 0 68172 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_741
timestamp 1644511149
transform 1 0 69276 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_753
timestamp 1644511149
transform 1 0 70380 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_765
timestamp 1644511149
transform 1 0 71484 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_777
timestamp 1644511149
transform 1 0 72588 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_783
timestamp 1644511149
transform 1 0 73140 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_785
timestamp 1644511149
transform 1 0 73324 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_797
timestamp 1644511149
transform 1 0 74428 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_809
timestamp 1644511149
transform 1 0 75532 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_821
timestamp 1644511149
transform 1 0 76636 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_833
timestamp 1644511149
transform 1 0 77740 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_839
timestamp 1644511149
transform 1 0 78292 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_841
timestamp 1644511149
transform 1 0 78476 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_3
timestamp 1644511149
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_15
timestamp 1644511149
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1644511149
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_29
timestamp 1644511149
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_41
timestamp 1644511149
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_53
timestamp 1644511149
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_65
timestamp 1644511149
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 1644511149
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1644511149
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_85
timestamp 1644511149
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_97
timestamp 1644511149
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_109
timestamp 1644511149
transform 1 0 11132 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_121
timestamp 1644511149
transform 1 0 12236 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_133
timestamp 1644511149
transform 1 0 13340 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 1644511149
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_141
timestamp 1644511149
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_153
timestamp 1644511149
transform 1 0 15180 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_165
timestamp 1644511149
transform 1 0 16284 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_177
timestamp 1644511149
transform 1 0 17388 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_189
timestamp 1644511149
transform 1 0 18492 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_195
timestamp 1644511149
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_197
timestamp 1644511149
transform 1 0 19228 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_209
timestamp 1644511149
transform 1 0 20332 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_221
timestamp 1644511149
transform 1 0 21436 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_233
timestamp 1644511149
transform 1 0 22540 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_245
timestamp 1644511149
transform 1 0 23644 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_251
timestamp 1644511149
transform 1 0 24196 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_253
timestamp 1644511149
transform 1 0 24380 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_265
timestamp 1644511149
transform 1 0 25484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_277
timestamp 1644511149
transform 1 0 26588 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_289
timestamp 1644511149
transform 1 0 27692 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_301
timestamp 1644511149
transform 1 0 28796 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_307
timestamp 1644511149
transform 1 0 29348 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_309
timestamp 1644511149
transform 1 0 29532 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_321
timestamp 1644511149
transform 1 0 30636 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_333
timestamp 1644511149
transform 1 0 31740 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_345
timestamp 1644511149
transform 1 0 32844 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_357
timestamp 1644511149
transform 1 0 33948 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_363
timestamp 1644511149
transform 1 0 34500 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_365
timestamp 1644511149
transform 1 0 34684 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_377
timestamp 1644511149
transform 1 0 35788 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_389
timestamp 1644511149
transform 1 0 36892 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_401
timestamp 1644511149
transform 1 0 37996 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_413
timestamp 1644511149
transform 1 0 39100 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_419
timestamp 1644511149
transform 1 0 39652 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_421
timestamp 1644511149
transform 1 0 39836 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_433
timestamp 1644511149
transform 1 0 40940 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_445
timestamp 1644511149
transform 1 0 42044 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_457
timestamp 1644511149
transform 1 0 43148 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_469
timestamp 1644511149
transform 1 0 44252 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_475
timestamp 1644511149
transform 1 0 44804 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_477
timestamp 1644511149
transform 1 0 44988 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_489
timestamp 1644511149
transform 1 0 46092 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_501
timestamp 1644511149
transform 1 0 47196 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_513
timestamp 1644511149
transform 1 0 48300 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_525
timestamp 1644511149
transform 1 0 49404 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_531
timestamp 1644511149
transform 1 0 49956 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_533
timestamp 1644511149
transform 1 0 50140 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_545
timestamp 1644511149
transform 1 0 51244 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_557
timestamp 1644511149
transform 1 0 52348 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_569
timestamp 1644511149
transform 1 0 53452 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_581
timestamp 1644511149
transform 1 0 54556 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_587
timestamp 1644511149
transform 1 0 55108 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_589
timestamp 1644511149
transform 1 0 55292 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_601
timestamp 1644511149
transform 1 0 56396 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_613
timestamp 1644511149
transform 1 0 57500 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_625
timestamp 1644511149
transform 1 0 58604 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_637
timestamp 1644511149
transform 1 0 59708 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_643
timestamp 1644511149
transform 1 0 60260 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_645
timestamp 1644511149
transform 1 0 60444 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_657
timestamp 1644511149
transform 1 0 61548 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_669
timestamp 1644511149
transform 1 0 62652 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_681
timestamp 1644511149
transform 1 0 63756 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_693
timestamp 1644511149
transform 1 0 64860 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_699
timestamp 1644511149
transform 1 0 65412 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_701
timestamp 1644511149
transform 1 0 65596 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_713
timestamp 1644511149
transform 1 0 66700 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_725
timestamp 1644511149
transform 1 0 67804 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_737
timestamp 1644511149
transform 1 0 68908 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_749
timestamp 1644511149
transform 1 0 70012 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_755
timestamp 1644511149
transform 1 0 70564 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_757
timestamp 1644511149
transform 1 0 70748 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_769
timestamp 1644511149
transform 1 0 71852 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_781
timestamp 1644511149
transform 1 0 72956 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_793
timestamp 1644511149
transform 1 0 74060 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_805
timestamp 1644511149
transform 1 0 75164 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_811
timestamp 1644511149
transform 1 0 75716 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_813
timestamp 1644511149
transform 1 0 75900 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_825
timestamp 1644511149
transform 1 0 77004 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_837
timestamp 1644511149
transform 1 0 78108 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_841
timestamp 1644511149
transform 1 0 78476 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_9
timestamp 1644511149
transform 1 0 1932 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_21
timestamp 1644511149
transform 1 0 3036 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_33
timestamp 1644511149
transform 1 0 4140 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_45
timestamp 1644511149
transform 1 0 5244 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_53
timestamp 1644511149
transform 1 0 5980 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_57
timestamp 1644511149
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_69
timestamp 1644511149
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_81
timestamp 1644511149
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_93
timestamp 1644511149
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_105
timestamp 1644511149
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1644511149
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_113
timestamp 1644511149
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_125
timestamp 1644511149
transform 1 0 12604 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_137
timestamp 1644511149
transform 1 0 13708 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_149
timestamp 1644511149
transform 1 0 14812 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_161
timestamp 1644511149
transform 1 0 15916 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_167
timestamp 1644511149
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_169
timestamp 1644511149
transform 1 0 16652 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_181
timestamp 1644511149
transform 1 0 17756 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_193
timestamp 1644511149
transform 1 0 18860 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_205
timestamp 1644511149
transform 1 0 19964 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_217
timestamp 1644511149
transform 1 0 21068 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_223
timestamp 1644511149
transform 1 0 21620 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_225
timestamp 1644511149
transform 1 0 21804 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_237
timestamp 1644511149
transform 1 0 22908 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_249
timestamp 1644511149
transform 1 0 24012 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_261
timestamp 1644511149
transform 1 0 25116 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_273
timestamp 1644511149
transform 1 0 26220 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_279
timestamp 1644511149
transform 1 0 26772 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_281
timestamp 1644511149
transform 1 0 26956 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_293
timestamp 1644511149
transform 1 0 28060 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_305
timestamp 1644511149
transform 1 0 29164 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_317
timestamp 1644511149
transform 1 0 30268 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_329
timestamp 1644511149
transform 1 0 31372 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_335
timestamp 1644511149
transform 1 0 31924 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_337
timestamp 1644511149
transform 1 0 32108 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_349
timestamp 1644511149
transform 1 0 33212 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_361
timestamp 1644511149
transform 1 0 34316 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_373
timestamp 1644511149
transform 1 0 35420 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_385
timestamp 1644511149
transform 1 0 36524 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_391
timestamp 1644511149
transform 1 0 37076 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_393
timestamp 1644511149
transform 1 0 37260 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_405
timestamp 1644511149
transform 1 0 38364 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_417
timestamp 1644511149
transform 1 0 39468 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_429
timestamp 1644511149
transform 1 0 40572 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_441
timestamp 1644511149
transform 1 0 41676 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_447
timestamp 1644511149
transform 1 0 42228 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_449
timestamp 1644511149
transform 1 0 42412 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_461
timestamp 1644511149
transform 1 0 43516 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_473
timestamp 1644511149
transform 1 0 44620 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_485
timestamp 1644511149
transform 1 0 45724 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_497
timestamp 1644511149
transform 1 0 46828 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_503
timestamp 1644511149
transform 1 0 47380 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_505
timestamp 1644511149
transform 1 0 47564 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_517
timestamp 1644511149
transform 1 0 48668 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_529
timestamp 1644511149
transform 1 0 49772 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_541
timestamp 1644511149
transform 1 0 50876 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_553
timestamp 1644511149
transform 1 0 51980 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_559
timestamp 1644511149
transform 1 0 52532 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_561
timestamp 1644511149
transform 1 0 52716 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_573
timestamp 1644511149
transform 1 0 53820 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_585
timestamp 1644511149
transform 1 0 54924 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_597
timestamp 1644511149
transform 1 0 56028 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_609
timestamp 1644511149
transform 1 0 57132 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_615
timestamp 1644511149
transform 1 0 57684 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_617
timestamp 1644511149
transform 1 0 57868 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_629
timestamp 1644511149
transform 1 0 58972 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_641
timestamp 1644511149
transform 1 0 60076 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_653
timestamp 1644511149
transform 1 0 61180 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_665
timestamp 1644511149
transform 1 0 62284 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_671
timestamp 1644511149
transform 1 0 62836 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_673
timestamp 1644511149
transform 1 0 63020 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_685
timestamp 1644511149
transform 1 0 64124 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_697
timestamp 1644511149
transform 1 0 65228 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_709
timestamp 1644511149
transform 1 0 66332 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_721
timestamp 1644511149
transform 1 0 67436 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_727
timestamp 1644511149
transform 1 0 67988 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_729
timestamp 1644511149
transform 1 0 68172 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_741
timestamp 1644511149
transform 1 0 69276 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_753
timestamp 1644511149
transform 1 0 70380 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_765
timestamp 1644511149
transform 1 0 71484 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_777
timestamp 1644511149
transform 1 0 72588 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_783
timestamp 1644511149
transform 1 0 73140 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_785
timestamp 1644511149
transform 1 0 73324 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_797
timestamp 1644511149
transform 1 0 74428 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_809
timestamp 1644511149
transform 1 0 75532 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_821
timestamp 1644511149
transform 1 0 76636 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_833
timestamp 1644511149
transform 1 0 77740 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_839
timestamp 1644511149
transform 1 0 78292 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_841
timestamp 1644511149
transform 1 0 78476 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_3
timestamp 1644511149
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_15
timestamp 1644511149
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1644511149
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_29
timestamp 1644511149
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_41
timestamp 1644511149
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_53
timestamp 1644511149
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_65
timestamp 1644511149
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_77
timestamp 1644511149
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1644511149
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_85
timestamp 1644511149
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_97
timestamp 1644511149
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_109
timestamp 1644511149
transform 1 0 11132 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_121
timestamp 1644511149
transform 1 0 12236 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_133
timestamp 1644511149
transform 1 0 13340 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_139
timestamp 1644511149
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_141
timestamp 1644511149
transform 1 0 14076 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_153
timestamp 1644511149
transform 1 0 15180 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_165
timestamp 1644511149
transform 1 0 16284 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_177
timestamp 1644511149
transform 1 0 17388 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_189
timestamp 1644511149
transform 1 0 18492 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_195
timestamp 1644511149
transform 1 0 19044 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_197
timestamp 1644511149
transform 1 0 19228 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_209
timestamp 1644511149
transform 1 0 20332 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_221
timestamp 1644511149
transform 1 0 21436 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_233
timestamp 1644511149
transform 1 0 22540 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_245
timestamp 1644511149
transform 1 0 23644 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_251
timestamp 1644511149
transform 1 0 24196 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_253
timestamp 1644511149
transform 1 0 24380 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_265
timestamp 1644511149
transform 1 0 25484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_277
timestamp 1644511149
transform 1 0 26588 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_289
timestamp 1644511149
transform 1 0 27692 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_301
timestamp 1644511149
transform 1 0 28796 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_307
timestamp 1644511149
transform 1 0 29348 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_309
timestamp 1644511149
transform 1 0 29532 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_321
timestamp 1644511149
transform 1 0 30636 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_333
timestamp 1644511149
transform 1 0 31740 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_345
timestamp 1644511149
transform 1 0 32844 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_357
timestamp 1644511149
transform 1 0 33948 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_363
timestamp 1644511149
transform 1 0 34500 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_365
timestamp 1644511149
transform 1 0 34684 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_377
timestamp 1644511149
transform 1 0 35788 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_389
timestamp 1644511149
transform 1 0 36892 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_401
timestamp 1644511149
transform 1 0 37996 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_413
timestamp 1644511149
transform 1 0 39100 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_419
timestamp 1644511149
transform 1 0 39652 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_421
timestamp 1644511149
transform 1 0 39836 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_18_431
timestamp 1644511149
transform 1 0 40756 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_443
timestamp 1644511149
transform 1 0 41860 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_455
timestamp 1644511149
transform 1 0 42964 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_467
timestamp 1644511149
transform 1 0 44068 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_475
timestamp 1644511149
transform 1 0 44804 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_477
timestamp 1644511149
transform 1 0 44988 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_489
timestamp 1644511149
transform 1 0 46092 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_501
timestamp 1644511149
transform 1 0 47196 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_513
timestamp 1644511149
transform 1 0 48300 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_525
timestamp 1644511149
transform 1 0 49404 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_531
timestamp 1644511149
transform 1 0 49956 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_533
timestamp 1644511149
transform 1 0 50140 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_545
timestamp 1644511149
transform 1 0 51244 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_557
timestamp 1644511149
transform 1 0 52348 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_569
timestamp 1644511149
transform 1 0 53452 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_581
timestamp 1644511149
transform 1 0 54556 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_587
timestamp 1644511149
transform 1 0 55108 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_589
timestamp 1644511149
transform 1 0 55292 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_601
timestamp 1644511149
transform 1 0 56396 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_613
timestamp 1644511149
transform 1 0 57500 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_625
timestamp 1644511149
transform 1 0 58604 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_637
timestamp 1644511149
transform 1 0 59708 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_643
timestamp 1644511149
transform 1 0 60260 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_645
timestamp 1644511149
transform 1 0 60444 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_657
timestamp 1644511149
transform 1 0 61548 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_669
timestamp 1644511149
transform 1 0 62652 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_681
timestamp 1644511149
transform 1 0 63756 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_693
timestamp 1644511149
transform 1 0 64860 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_699
timestamp 1644511149
transform 1 0 65412 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_701
timestamp 1644511149
transform 1 0 65596 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_713
timestamp 1644511149
transform 1 0 66700 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_725
timestamp 1644511149
transform 1 0 67804 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_737
timestamp 1644511149
transform 1 0 68908 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_749
timestamp 1644511149
transform 1 0 70012 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_755
timestamp 1644511149
transform 1 0 70564 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_757
timestamp 1644511149
transform 1 0 70748 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_769
timestamp 1644511149
transform 1 0 71852 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_781
timestamp 1644511149
transform 1 0 72956 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_793
timestamp 1644511149
transform 1 0 74060 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_805
timestamp 1644511149
transform 1 0 75164 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_811
timestamp 1644511149
transform 1 0 75716 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_813
timestamp 1644511149
transform 1 0 75900 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_825
timestamp 1644511149
transform 1 0 77004 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_837
timestamp 1644511149
transform 1 0 78108 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_841
timestamp 1644511149
transform 1 0 78476 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_3
timestamp 1644511149
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_15
timestamp 1644511149
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_27
timestamp 1644511149
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_39
timestamp 1644511149
transform 1 0 4692 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_51
timestamp 1644511149
transform 1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1644511149
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_57
timestamp 1644511149
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_69
timestamp 1644511149
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_81
timestamp 1644511149
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_93
timestamp 1644511149
transform 1 0 9660 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_105
timestamp 1644511149
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1644511149
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_113
timestamp 1644511149
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_125
timestamp 1644511149
transform 1 0 12604 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_137
timestamp 1644511149
transform 1 0 13708 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_149
timestamp 1644511149
transform 1 0 14812 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_161
timestamp 1644511149
transform 1 0 15916 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_167
timestamp 1644511149
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_169
timestamp 1644511149
transform 1 0 16652 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_181
timestamp 1644511149
transform 1 0 17756 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_193
timestamp 1644511149
transform 1 0 18860 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_205
timestamp 1644511149
transform 1 0 19964 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_217
timestamp 1644511149
transform 1 0 21068 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_223
timestamp 1644511149
transform 1 0 21620 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_225
timestamp 1644511149
transform 1 0 21804 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_237
timestamp 1644511149
transform 1 0 22908 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_249
timestamp 1644511149
transform 1 0 24012 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_261
timestamp 1644511149
transform 1 0 25116 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_273
timestamp 1644511149
transform 1 0 26220 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_279
timestamp 1644511149
transform 1 0 26772 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_281
timestamp 1644511149
transform 1 0 26956 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_293
timestamp 1644511149
transform 1 0 28060 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_305
timestamp 1644511149
transform 1 0 29164 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_317
timestamp 1644511149
transform 1 0 30268 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_329
timestamp 1644511149
transform 1 0 31372 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_335
timestamp 1644511149
transform 1 0 31924 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_337
timestamp 1644511149
transform 1 0 32108 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_349
timestamp 1644511149
transform 1 0 33212 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_361
timestamp 1644511149
transform 1 0 34316 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_373
timestamp 1644511149
transform 1 0 35420 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_385
timestamp 1644511149
transform 1 0 36524 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_391
timestamp 1644511149
transform 1 0 37076 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_393
timestamp 1644511149
transform 1 0 37260 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_405
timestamp 1644511149
transform 1 0 38364 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_417
timestamp 1644511149
transform 1 0 39468 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_429
timestamp 1644511149
transform 1 0 40572 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_441
timestamp 1644511149
transform 1 0 41676 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_447
timestamp 1644511149
transform 1 0 42228 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_449
timestamp 1644511149
transform 1 0 42412 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_461
timestamp 1644511149
transform 1 0 43516 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_473
timestamp 1644511149
transform 1 0 44620 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_485
timestamp 1644511149
transform 1 0 45724 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_497
timestamp 1644511149
transform 1 0 46828 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_503
timestamp 1644511149
transform 1 0 47380 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_505
timestamp 1644511149
transform 1 0 47564 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_517
timestamp 1644511149
transform 1 0 48668 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_529
timestamp 1644511149
transform 1 0 49772 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_541
timestamp 1644511149
transform 1 0 50876 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_553
timestamp 1644511149
transform 1 0 51980 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_559
timestamp 1644511149
transform 1 0 52532 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_561
timestamp 1644511149
transform 1 0 52716 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_573
timestamp 1644511149
transform 1 0 53820 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_585
timestamp 1644511149
transform 1 0 54924 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_597
timestamp 1644511149
transform 1 0 56028 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_609
timestamp 1644511149
transform 1 0 57132 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_615
timestamp 1644511149
transform 1 0 57684 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_617
timestamp 1644511149
transform 1 0 57868 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_629
timestamp 1644511149
transform 1 0 58972 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_641
timestamp 1644511149
transform 1 0 60076 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_653
timestamp 1644511149
transform 1 0 61180 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_665
timestamp 1644511149
transform 1 0 62284 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_671
timestamp 1644511149
transform 1 0 62836 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_673
timestamp 1644511149
transform 1 0 63020 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_685
timestamp 1644511149
transform 1 0 64124 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_697
timestamp 1644511149
transform 1 0 65228 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_709
timestamp 1644511149
transform 1 0 66332 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_721
timestamp 1644511149
transform 1 0 67436 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_727
timestamp 1644511149
transform 1 0 67988 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_729
timestamp 1644511149
transform 1 0 68172 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_741
timestamp 1644511149
transform 1 0 69276 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_753
timestamp 1644511149
transform 1 0 70380 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_765
timestamp 1644511149
transform 1 0 71484 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_777
timestamp 1644511149
transform 1 0 72588 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_783
timestamp 1644511149
transform 1 0 73140 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_785
timestamp 1644511149
transform 1 0 73324 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_797
timestamp 1644511149
transform 1 0 74428 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_809
timestamp 1644511149
transform 1 0 75532 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_821
timestamp 1644511149
transform 1 0 76636 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_829
timestamp 1644511149
transform 1 0 77372 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_836
timestamp 1644511149
transform 1 0 78016 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_841
timestamp 1644511149
transform 1 0 78476 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_3
timestamp 1644511149
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_15
timestamp 1644511149
transform 1 0 2484 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_20_21
timestamp 1644511149
transform 1 0 3036 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1644511149
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_29
timestamp 1644511149
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_41
timestamp 1644511149
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_53
timestamp 1644511149
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_65
timestamp 1644511149
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_77
timestamp 1644511149
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1644511149
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_85
timestamp 1644511149
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_97
timestamp 1644511149
transform 1 0 10028 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_109
timestamp 1644511149
transform 1 0 11132 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_121
timestamp 1644511149
transform 1 0 12236 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_133
timestamp 1644511149
transform 1 0 13340 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp 1644511149
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_141
timestamp 1644511149
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_153
timestamp 1644511149
transform 1 0 15180 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_165
timestamp 1644511149
transform 1 0 16284 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_177
timestamp 1644511149
transform 1 0 17388 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_189
timestamp 1644511149
transform 1 0 18492 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_195
timestamp 1644511149
transform 1 0 19044 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_197
timestamp 1644511149
transform 1 0 19228 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_209
timestamp 1644511149
transform 1 0 20332 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_221
timestamp 1644511149
transform 1 0 21436 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_233
timestamp 1644511149
transform 1 0 22540 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_245
timestamp 1644511149
transform 1 0 23644 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_251
timestamp 1644511149
transform 1 0 24196 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_253
timestamp 1644511149
transform 1 0 24380 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_265
timestamp 1644511149
transform 1 0 25484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_277
timestamp 1644511149
transform 1 0 26588 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_289
timestamp 1644511149
transform 1 0 27692 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_301
timestamp 1644511149
transform 1 0 28796 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_307
timestamp 1644511149
transform 1 0 29348 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_309
timestamp 1644511149
transform 1 0 29532 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_321
timestamp 1644511149
transform 1 0 30636 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_333
timestamp 1644511149
transform 1 0 31740 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_345
timestamp 1644511149
transform 1 0 32844 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_357
timestamp 1644511149
transform 1 0 33948 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_363
timestamp 1644511149
transform 1 0 34500 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_365
timestamp 1644511149
transform 1 0 34684 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_377
timestamp 1644511149
transform 1 0 35788 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_389
timestamp 1644511149
transform 1 0 36892 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_401
timestamp 1644511149
transform 1 0 37996 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_413
timestamp 1644511149
transform 1 0 39100 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_419
timestamp 1644511149
transform 1 0 39652 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_421
timestamp 1644511149
transform 1 0 39836 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_433
timestamp 1644511149
transform 1 0 40940 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_445
timestamp 1644511149
transform 1 0 42044 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_457
timestamp 1644511149
transform 1 0 43148 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_469
timestamp 1644511149
transform 1 0 44252 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_475
timestamp 1644511149
transform 1 0 44804 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_477
timestamp 1644511149
transform 1 0 44988 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_489
timestamp 1644511149
transform 1 0 46092 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_501
timestamp 1644511149
transform 1 0 47196 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_513
timestamp 1644511149
transform 1 0 48300 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_525
timestamp 1644511149
transform 1 0 49404 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_531
timestamp 1644511149
transform 1 0 49956 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_533
timestamp 1644511149
transform 1 0 50140 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_545
timestamp 1644511149
transform 1 0 51244 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_557
timestamp 1644511149
transform 1 0 52348 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_569
timestamp 1644511149
transform 1 0 53452 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_581
timestamp 1644511149
transform 1 0 54556 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_587
timestamp 1644511149
transform 1 0 55108 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_589
timestamp 1644511149
transform 1 0 55292 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_601
timestamp 1644511149
transform 1 0 56396 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_613
timestamp 1644511149
transform 1 0 57500 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_625
timestamp 1644511149
transform 1 0 58604 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_637
timestamp 1644511149
transform 1 0 59708 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_643
timestamp 1644511149
transform 1 0 60260 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_645
timestamp 1644511149
transform 1 0 60444 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_657
timestamp 1644511149
transform 1 0 61548 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_669
timestamp 1644511149
transform 1 0 62652 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_681
timestamp 1644511149
transform 1 0 63756 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_693
timestamp 1644511149
transform 1 0 64860 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_699
timestamp 1644511149
transform 1 0 65412 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_701
timestamp 1644511149
transform 1 0 65596 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_713
timestamp 1644511149
transform 1 0 66700 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_725
timestamp 1644511149
transform 1 0 67804 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_737
timestamp 1644511149
transform 1 0 68908 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_749
timestamp 1644511149
transform 1 0 70012 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_755
timestamp 1644511149
transform 1 0 70564 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_757
timestamp 1644511149
transform 1 0 70748 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_769
timestamp 1644511149
transform 1 0 71852 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_781
timestamp 1644511149
transform 1 0 72956 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_793
timestamp 1644511149
transform 1 0 74060 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_805
timestamp 1644511149
transform 1 0 75164 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_811
timestamp 1644511149
transform 1 0 75716 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_813
timestamp 1644511149
transform 1 0 75900 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_825
timestamp 1644511149
transform 1 0 77004 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_837
timestamp 1644511149
transform 1 0 78108 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_841
timestamp 1644511149
transform 1 0 78476 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_3
timestamp 1644511149
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_15
timestamp 1644511149
transform 1 0 2484 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_27
timestamp 1644511149
transform 1 0 3588 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_39
timestamp 1644511149
transform 1 0 4692 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_51
timestamp 1644511149
transform 1 0 5796 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1644511149
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_57
timestamp 1644511149
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_69
timestamp 1644511149
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_81
timestamp 1644511149
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_93
timestamp 1644511149
transform 1 0 9660 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_105
timestamp 1644511149
transform 1 0 10764 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1644511149
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_113
timestamp 1644511149
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_125
timestamp 1644511149
transform 1 0 12604 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_137
timestamp 1644511149
transform 1 0 13708 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_149
timestamp 1644511149
transform 1 0 14812 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_161
timestamp 1644511149
transform 1 0 15916 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_167
timestamp 1644511149
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_169
timestamp 1644511149
transform 1 0 16652 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_181
timestamp 1644511149
transform 1 0 17756 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_193
timestamp 1644511149
transform 1 0 18860 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_205
timestamp 1644511149
transform 1 0 19964 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_217
timestamp 1644511149
transform 1 0 21068 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_223
timestamp 1644511149
transform 1 0 21620 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_225
timestamp 1644511149
transform 1 0 21804 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_237
timestamp 1644511149
transform 1 0 22908 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_249
timestamp 1644511149
transform 1 0 24012 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_261
timestamp 1644511149
transform 1 0 25116 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_273
timestamp 1644511149
transform 1 0 26220 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_279
timestamp 1644511149
transform 1 0 26772 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_281
timestamp 1644511149
transform 1 0 26956 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_293
timestamp 1644511149
transform 1 0 28060 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_305
timestamp 1644511149
transform 1 0 29164 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_317
timestamp 1644511149
transform 1 0 30268 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_329
timestamp 1644511149
transform 1 0 31372 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_335
timestamp 1644511149
transform 1 0 31924 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_337
timestamp 1644511149
transform 1 0 32108 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_349
timestamp 1644511149
transform 1 0 33212 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_361
timestamp 1644511149
transform 1 0 34316 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_373
timestamp 1644511149
transform 1 0 35420 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_385
timestamp 1644511149
transform 1 0 36524 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_391
timestamp 1644511149
transform 1 0 37076 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_393
timestamp 1644511149
transform 1 0 37260 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_405
timestamp 1644511149
transform 1 0 38364 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_417
timestamp 1644511149
transform 1 0 39468 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_429
timestamp 1644511149
transform 1 0 40572 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_441
timestamp 1644511149
transform 1 0 41676 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_447
timestamp 1644511149
transform 1 0 42228 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_449
timestamp 1644511149
transform 1 0 42412 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_461
timestamp 1644511149
transform 1 0 43516 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_473
timestamp 1644511149
transform 1 0 44620 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_485
timestamp 1644511149
transform 1 0 45724 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_497
timestamp 1644511149
transform 1 0 46828 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_503
timestamp 1644511149
transform 1 0 47380 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_505
timestamp 1644511149
transform 1 0 47564 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_517
timestamp 1644511149
transform 1 0 48668 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_529
timestamp 1644511149
transform 1 0 49772 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_541
timestamp 1644511149
transform 1 0 50876 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_553
timestamp 1644511149
transform 1 0 51980 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_559
timestamp 1644511149
transform 1 0 52532 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_561
timestamp 1644511149
transform 1 0 52716 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_573
timestamp 1644511149
transform 1 0 53820 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_585
timestamp 1644511149
transform 1 0 54924 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_597
timestamp 1644511149
transform 1 0 56028 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_609
timestamp 1644511149
transform 1 0 57132 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_615
timestamp 1644511149
transform 1 0 57684 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_617
timestamp 1644511149
transform 1 0 57868 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_629
timestamp 1644511149
transform 1 0 58972 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_641
timestamp 1644511149
transform 1 0 60076 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_653
timestamp 1644511149
transform 1 0 61180 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_665
timestamp 1644511149
transform 1 0 62284 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_671
timestamp 1644511149
transform 1 0 62836 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_673
timestamp 1644511149
transform 1 0 63020 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_685
timestamp 1644511149
transform 1 0 64124 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_697
timestamp 1644511149
transform 1 0 65228 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_709
timestamp 1644511149
transform 1 0 66332 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_721
timestamp 1644511149
transform 1 0 67436 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_727
timestamp 1644511149
transform 1 0 67988 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_729
timestamp 1644511149
transform 1 0 68172 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_741
timestamp 1644511149
transform 1 0 69276 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_753
timestamp 1644511149
transform 1 0 70380 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_765
timestamp 1644511149
transform 1 0 71484 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_777
timestamp 1644511149
transform 1 0 72588 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_783
timestamp 1644511149
transform 1 0 73140 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_785
timestamp 1644511149
transform 1 0 73324 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_797
timestamp 1644511149
transform 1 0 74428 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_809
timestamp 1644511149
transform 1 0 75532 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_821
timestamp 1644511149
transform 1 0 76636 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_833
timestamp 1644511149
transform 1 0 77740 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_839
timestamp 1644511149
transform 1 0 78292 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_841
timestamp 1644511149
transform 1 0 78476 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_3
timestamp 1644511149
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_15
timestamp 1644511149
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1644511149
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_29
timestamp 1644511149
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_41
timestamp 1644511149
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_53
timestamp 1644511149
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_65
timestamp 1644511149
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_77
timestamp 1644511149
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1644511149
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_85
timestamp 1644511149
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_97
timestamp 1644511149
transform 1 0 10028 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_109
timestamp 1644511149
transform 1 0 11132 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_121
timestamp 1644511149
transform 1 0 12236 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_133
timestamp 1644511149
transform 1 0 13340 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_139
timestamp 1644511149
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_141
timestamp 1644511149
transform 1 0 14076 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_153
timestamp 1644511149
transform 1 0 15180 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_165
timestamp 1644511149
transform 1 0 16284 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_177
timestamp 1644511149
transform 1 0 17388 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_189
timestamp 1644511149
transform 1 0 18492 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_195
timestamp 1644511149
transform 1 0 19044 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_197
timestamp 1644511149
transform 1 0 19228 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_209
timestamp 1644511149
transform 1 0 20332 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_221
timestamp 1644511149
transform 1 0 21436 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_233
timestamp 1644511149
transform 1 0 22540 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_245
timestamp 1644511149
transform 1 0 23644 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_251
timestamp 1644511149
transform 1 0 24196 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_253
timestamp 1644511149
transform 1 0 24380 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_265
timestamp 1644511149
transform 1 0 25484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_277
timestamp 1644511149
transform 1 0 26588 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_289
timestamp 1644511149
transform 1 0 27692 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_301
timestamp 1644511149
transform 1 0 28796 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_307
timestamp 1644511149
transform 1 0 29348 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_309
timestamp 1644511149
transform 1 0 29532 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_321
timestamp 1644511149
transform 1 0 30636 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_333
timestamp 1644511149
transform 1 0 31740 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_345
timestamp 1644511149
transform 1 0 32844 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_357
timestamp 1644511149
transform 1 0 33948 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_363
timestamp 1644511149
transform 1 0 34500 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_365
timestamp 1644511149
transform 1 0 34684 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_377
timestamp 1644511149
transform 1 0 35788 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_389
timestamp 1644511149
transform 1 0 36892 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_401
timestamp 1644511149
transform 1 0 37996 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_413
timestamp 1644511149
transform 1 0 39100 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_419
timestamp 1644511149
transform 1 0 39652 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_421
timestamp 1644511149
transform 1 0 39836 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_433
timestamp 1644511149
transform 1 0 40940 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_445
timestamp 1644511149
transform 1 0 42044 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_457
timestamp 1644511149
transform 1 0 43148 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_469
timestamp 1644511149
transform 1 0 44252 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_475
timestamp 1644511149
transform 1 0 44804 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_477
timestamp 1644511149
transform 1 0 44988 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_489
timestamp 1644511149
transform 1 0 46092 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_501
timestamp 1644511149
transform 1 0 47196 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_513
timestamp 1644511149
transform 1 0 48300 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_525
timestamp 1644511149
transform 1 0 49404 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_531
timestamp 1644511149
transform 1 0 49956 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_533
timestamp 1644511149
transform 1 0 50140 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_545
timestamp 1644511149
transform 1 0 51244 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_557
timestamp 1644511149
transform 1 0 52348 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_569
timestamp 1644511149
transform 1 0 53452 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_581
timestamp 1644511149
transform 1 0 54556 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_587
timestamp 1644511149
transform 1 0 55108 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_589
timestamp 1644511149
transform 1 0 55292 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_601
timestamp 1644511149
transform 1 0 56396 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_613
timestamp 1644511149
transform 1 0 57500 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_625
timestamp 1644511149
transform 1 0 58604 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_637
timestamp 1644511149
transform 1 0 59708 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_643
timestamp 1644511149
transform 1 0 60260 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_645
timestamp 1644511149
transform 1 0 60444 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_657
timestamp 1644511149
transform 1 0 61548 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_669
timestamp 1644511149
transform 1 0 62652 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_681
timestamp 1644511149
transform 1 0 63756 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_693
timestamp 1644511149
transform 1 0 64860 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_699
timestamp 1644511149
transform 1 0 65412 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_701
timestamp 1644511149
transform 1 0 65596 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_713
timestamp 1644511149
transform 1 0 66700 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_725
timestamp 1644511149
transform 1 0 67804 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_737
timestamp 1644511149
transform 1 0 68908 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_749
timestamp 1644511149
transform 1 0 70012 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_755
timestamp 1644511149
transform 1 0 70564 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_757
timestamp 1644511149
transform 1 0 70748 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_769
timestamp 1644511149
transform 1 0 71852 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_781
timestamp 1644511149
transform 1 0 72956 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_793
timestamp 1644511149
transform 1 0 74060 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_805
timestamp 1644511149
transform 1 0 75164 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_811
timestamp 1644511149
transform 1 0 75716 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_813
timestamp 1644511149
transform 1 0 75900 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_825
timestamp 1644511149
transform 1 0 77004 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_837
timestamp 1644511149
transform 1 0 78108 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_841
timestamp 1644511149
transform 1 0 78476 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_3
timestamp 1644511149
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_15
timestamp 1644511149
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_27
timestamp 1644511149
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_39
timestamp 1644511149
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_51
timestamp 1644511149
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1644511149
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_57
timestamp 1644511149
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_69
timestamp 1644511149
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_81
timestamp 1644511149
transform 1 0 8556 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_93
timestamp 1644511149
transform 1 0 9660 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_105
timestamp 1644511149
transform 1 0 10764 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 1644511149
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_113
timestamp 1644511149
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_125
timestamp 1644511149
transform 1 0 12604 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_137
timestamp 1644511149
transform 1 0 13708 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_149
timestamp 1644511149
transform 1 0 14812 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_161
timestamp 1644511149
transform 1 0 15916 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_167
timestamp 1644511149
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_169
timestamp 1644511149
transform 1 0 16652 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_181
timestamp 1644511149
transform 1 0 17756 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_193
timestamp 1644511149
transform 1 0 18860 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_205
timestamp 1644511149
transform 1 0 19964 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_217
timestamp 1644511149
transform 1 0 21068 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_223
timestamp 1644511149
transform 1 0 21620 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_225
timestamp 1644511149
transform 1 0 21804 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_237
timestamp 1644511149
transform 1 0 22908 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_249
timestamp 1644511149
transform 1 0 24012 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_261
timestamp 1644511149
transform 1 0 25116 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_273
timestamp 1644511149
transform 1 0 26220 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_279
timestamp 1644511149
transform 1 0 26772 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_281
timestamp 1644511149
transform 1 0 26956 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_293
timestamp 1644511149
transform 1 0 28060 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_305
timestamp 1644511149
transform 1 0 29164 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_317
timestamp 1644511149
transform 1 0 30268 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_329
timestamp 1644511149
transform 1 0 31372 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_335
timestamp 1644511149
transform 1 0 31924 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_337
timestamp 1644511149
transform 1 0 32108 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_349
timestamp 1644511149
transform 1 0 33212 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_361
timestamp 1644511149
transform 1 0 34316 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_373
timestamp 1644511149
transform 1 0 35420 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_385
timestamp 1644511149
transform 1 0 36524 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_391
timestamp 1644511149
transform 1 0 37076 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_393
timestamp 1644511149
transform 1 0 37260 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_405
timestamp 1644511149
transform 1 0 38364 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_417
timestamp 1644511149
transform 1 0 39468 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_429
timestamp 1644511149
transform 1 0 40572 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_441
timestamp 1644511149
transform 1 0 41676 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_447
timestamp 1644511149
transform 1 0 42228 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_449
timestamp 1644511149
transform 1 0 42412 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_461
timestamp 1644511149
transform 1 0 43516 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_473
timestamp 1644511149
transform 1 0 44620 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_485
timestamp 1644511149
transform 1 0 45724 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_497
timestamp 1644511149
transform 1 0 46828 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_503
timestamp 1644511149
transform 1 0 47380 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_505
timestamp 1644511149
transform 1 0 47564 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_517
timestamp 1644511149
transform 1 0 48668 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_529
timestamp 1644511149
transform 1 0 49772 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_541
timestamp 1644511149
transform 1 0 50876 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_553
timestamp 1644511149
transform 1 0 51980 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_559
timestamp 1644511149
transform 1 0 52532 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_561
timestamp 1644511149
transform 1 0 52716 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_573
timestamp 1644511149
transform 1 0 53820 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_585
timestamp 1644511149
transform 1 0 54924 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_597
timestamp 1644511149
transform 1 0 56028 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_609
timestamp 1644511149
transform 1 0 57132 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_615
timestamp 1644511149
transform 1 0 57684 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_617
timestamp 1644511149
transform 1 0 57868 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_629
timestamp 1644511149
transform 1 0 58972 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_641
timestamp 1644511149
transform 1 0 60076 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_653
timestamp 1644511149
transform 1 0 61180 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_665
timestamp 1644511149
transform 1 0 62284 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_671
timestamp 1644511149
transform 1 0 62836 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_673
timestamp 1644511149
transform 1 0 63020 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_685
timestamp 1644511149
transform 1 0 64124 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_697
timestamp 1644511149
transform 1 0 65228 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_709
timestamp 1644511149
transform 1 0 66332 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_721
timestamp 1644511149
transform 1 0 67436 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_727
timestamp 1644511149
transform 1 0 67988 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_729
timestamp 1644511149
transform 1 0 68172 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_741
timestamp 1644511149
transform 1 0 69276 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_753
timestamp 1644511149
transform 1 0 70380 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_765
timestamp 1644511149
transform 1 0 71484 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_777
timestamp 1644511149
transform 1 0 72588 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_783
timestamp 1644511149
transform 1 0 73140 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_785
timestamp 1644511149
transform 1 0 73324 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_797
timestamp 1644511149
transform 1 0 74428 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_809
timestamp 1644511149
transform 1 0 75532 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_821
timestamp 1644511149
transform 1 0 76636 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_833
timestamp 1644511149
transform 1 0 77740 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_839
timestamp 1644511149
transform 1 0 78292 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_23_841
timestamp 1644511149
transform 1 0 78476 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_3
timestamp 1644511149
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_15
timestamp 1644511149
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1644511149
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_29
timestamp 1644511149
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_41
timestamp 1644511149
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_53
timestamp 1644511149
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_65
timestamp 1644511149
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_77
timestamp 1644511149
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1644511149
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_85
timestamp 1644511149
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_97
timestamp 1644511149
transform 1 0 10028 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_109
timestamp 1644511149
transform 1 0 11132 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_121
timestamp 1644511149
transform 1 0 12236 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_133
timestamp 1644511149
transform 1 0 13340 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp 1644511149
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_141
timestamp 1644511149
transform 1 0 14076 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_153
timestamp 1644511149
transform 1 0 15180 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_165
timestamp 1644511149
transform 1 0 16284 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_177
timestamp 1644511149
transform 1 0 17388 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_189
timestamp 1644511149
transform 1 0 18492 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_195
timestamp 1644511149
transform 1 0 19044 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_197
timestamp 1644511149
transform 1 0 19228 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_209
timestamp 1644511149
transform 1 0 20332 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_221
timestamp 1644511149
transform 1 0 21436 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_233
timestamp 1644511149
transform 1 0 22540 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_245
timestamp 1644511149
transform 1 0 23644 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_251
timestamp 1644511149
transform 1 0 24196 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_253
timestamp 1644511149
transform 1 0 24380 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_265
timestamp 1644511149
transform 1 0 25484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_277
timestamp 1644511149
transform 1 0 26588 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_289
timestamp 1644511149
transform 1 0 27692 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_301
timestamp 1644511149
transform 1 0 28796 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_307
timestamp 1644511149
transform 1 0 29348 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_309
timestamp 1644511149
transform 1 0 29532 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_321
timestamp 1644511149
transform 1 0 30636 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_333
timestamp 1644511149
transform 1 0 31740 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_345
timestamp 1644511149
transform 1 0 32844 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_357
timestamp 1644511149
transform 1 0 33948 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_363
timestamp 1644511149
transform 1 0 34500 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_365
timestamp 1644511149
transform 1 0 34684 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_377
timestamp 1644511149
transform 1 0 35788 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_389
timestamp 1644511149
transform 1 0 36892 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_401
timestamp 1644511149
transform 1 0 37996 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_413
timestamp 1644511149
transform 1 0 39100 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_419
timestamp 1644511149
transform 1 0 39652 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_421
timestamp 1644511149
transform 1 0 39836 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_433
timestamp 1644511149
transform 1 0 40940 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_445
timestamp 1644511149
transform 1 0 42044 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_457
timestamp 1644511149
transform 1 0 43148 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_469
timestamp 1644511149
transform 1 0 44252 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_475
timestamp 1644511149
transform 1 0 44804 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_477
timestamp 1644511149
transform 1 0 44988 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_489
timestamp 1644511149
transform 1 0 46092 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_501
timestamp 1644511149
transform 1 0 47196 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_513
timestamp 1644511149
transform 1 0 48300 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_525
timestamp 1644511149
transform 1 0 49404 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_531
timestamp 1644511149
transform 1 0 49956 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_533
timestamp 1644511149
transform 1 0 50140 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_545
timestamp 1644511149
transform 1 0 51244 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_557
timestamp 1644511149
transform 1 0 52348 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_569
timestamp 1644511149
transform 1 0 53452 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_581
timestamp 1644511149
transform 1 0 54556 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_587
timestamp 1644511149
transform 1 0 55108 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_589
timestamp 1644511149
transform 1 0 55292 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_601
timestamp 1644511149
transform 1 0 56396 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_613
timestamp 1644511149
transform 1 0 57500 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_625
timestamp 1644511149
transform 1 0 58604 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_637
timestamp 1644511149
transform 1 0 59708 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_643
timestamp 1644511149
transform 1 0 60260 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_645
timestamp 1644511149
transform 1 0 60444 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_657
timestamp 1644511149
transform 1 0 61548 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_669
timestamp 1644511149
transform 1 0 62652 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_681
timestamp 1644511149
transform 1 0 63756 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_693
timestamp 1644511149
transform 1 0 64860 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_699
timestamp 1644511149
transform 1 0 65412 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_701
timestamp 1644511149
transform 1 0 65596 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_713
timestamp 1644511149
transform 1 0 66700 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_725
timestamp 1644511149
transform 1 0 67804 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_737
timestamp 1644511149
transform 1 0 68908 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_749
timestamp 1644511149
transform 1 0 70012 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_755
timestamp 1644511149
transform 1 0 70564 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_757
timestamp 1644511149
transform 1 0 70748 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_769
timestamp 1644511149
transform 1 0 71852 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_781
timestamp 1644511149
transform 1 0 72956 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_793
timestamp 1644511149
transform 1 0 74060 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_805
timestamp 1644511149
transform 1 0 75164 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_811
timestamp 1644511149
transform 1 0 75716 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_813
timestamp 1644511149
transform 1 0 75900 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_825
timestamp 1644511149
transform 1 0 77004 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_837
timestamp 1644511149
transform 1 0 78108 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_841
timestamp 1644511149
transform 1 0 78476 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_7
timestamp 1644511149
transform 1 0 1748 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_25_11
timestamp 1644511149
transform 1 0 2116 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_23
timestamp 1644511149
transform 1 0 3220 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_35
timestamp 1644511149
transform 1 0 4324 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_47
timestamp 1644511149
transform 1 0 5428 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_55
timestamp 1644511149
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_57
timestamp 1644511149
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_69
timestamp 1644511149
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_81
timestamp 1644511149
transform 1 0 8556 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_93
timestamp 1644511149
transform 1 0 9660 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_105
timestamp 1644511149
transform 1 0 10764 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 1644511149
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_113
timestamp 1644511149
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_125
timestamp 1644511149
transform 1 0 12604 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_137
timestamp 1644511149
transform 1 0 13708 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_149
timestamp 1644511149
transform 1 0 14812 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_161
timestamp 1644511149
transform 1 0 15916 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_167
timestamp 1644511149
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_169
timestamp 1644511149
transform 1 0 16652 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_181
timestamp 1644511149
transform 1 0 17756 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_193
timestamp 1644511149
transform 1 0 18860 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_205
timestamp 1644511149
transform 1 0 19964 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_217
timestamp 1644511149
transform 1 0 21068 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_223
timestamp 1644511149
transform 1 0 21620 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_225
timestamp 1644511149
transform 1 0 21804 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_237
timestamp 1644511149
transform 1 0 22908 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_249
timestamp 1644511149
transform 1 0 24012 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_261
timestamp 1644511149
transform 1 0 25116 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_273
timestamp 1644511149
transform 1 0 26220 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_279
timestamp 1644511149
transform 1 0 26772 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_281
timestamp 1644511149
transform 1 0 26956 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_293
timestamp 1644511149
transform 1 0 28060 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_305
timestamp 1644511149
transform 1 0 29164 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_317
timestamp 1644511149
transform 1 0 30268 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_329
timestamp 1644511149
transform 1 0 31372 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_335
timestamp 1644511149
transform 1 0 31924 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_337
timestamp 1644511149
transform 1 0 32108 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_349
timestamp 1644511149
transform 1 0 33212 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_361
timestamp 1644511149
transform 1 0 34316 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_373
timestamp 1644511149
transform 1 0 35420 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_385
timestamp 1644511149
transform 1 0 36524 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_391
timestamp 1644511149
transform 1 0 37076 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_393
timestamp 1644511149
transform 1 0 37260 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_405
timestamp 1644511149
transform 1 0 38364 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_417
timestamp 1644511149
transform 1 0 39468 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_429
timestamp 1644511149
transform 1 0 40572 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_441
timestamp 1644511149
transform 1 0 41676 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_447
timestamp 1644511149
transform 1 0 42228 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_449
timestamp 1644511149
transform 1 0 42412 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_461
timestamp 1644511149
transform 1 0 43516 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_473
timestamp 1644511149
transform 1 0 44620 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_485
timestamp 1644511149
transform 1 0 45724 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_497
timestamp 1644511149
transform 1 0 46828 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_503
timestamp 1644511149
transform 1 0 47380 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_505
timestamp 1644511149
transform 1 0 47564 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_517
timestamp 1644511149
transform 1 0 48668 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_529
timestamp 1644511149
transform 1 0 49772 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_541
timestamp 1644511149
transform 1 0 50876 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_553
timestamp 1644511149
transform 1 0 51980 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_559
timestamp 1644511149
transform 1 0 52532 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_561
timestamp 1644511149
transform 1 0 52716 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_573
timestamp 1644511149
transform 1 0 53820 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_585
timestamp 1644511149
transform 1 0 54924 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_597
timestamp 1644511149
transform 1 0 56028 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_609
timestamp 1644511149
transform 1 0 57132 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_615
timestamp 1644511149
transform 1 0 57684 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_617
timestamp 1644511149
transform 1 0 57868 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_629
timestamp 1644511149
transform 1 0 58972 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_641
timestamp 1644511149
transform 1 0 60076 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_653
timestamp 1644511149
transform 1 0 61180 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_665
timestamp 1644511149
transform 1 0 62284 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_671
timestamp 1644511149
transform 1 0 62836 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_673
timestamp 1644511149
transform 1 0 63020 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_685
timestamp 1644511149
transform 1 0 64124 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_697
timestamp 1644511149
transform 1 0 65228 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_709
timestamp 1644511149
transform 1 0 66332 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_721
timestamp 1644511149
transform 1 0 67436 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_727
timestamp 1644511149
transform 1 0 67988 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_729
timestamp 1644511149
transform 1 0 68172 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_741
timestamp 1644511149
transform 1 0 69276 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_753
timestamp 1644511149
transform 1 0 70380 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_765
timestamp 1644511149
transform 1 0 71484 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_777
timestamp 1644511149
transform 1 0 72588 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_783
timestamp 1644511149
transform 1 0 73140 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_785
timestamp 1644511149
transform 1 0 73324 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_797
timestamp 1644511149
transform 1 0 74428 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_809
timestamp 1644511149
transform 1 0 75532 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_821
timestamp 1644511149
transform 1 0 76636 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_833
timestamp 1644511149
transform 1 0 77740 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_839
timestamp 1644511149
transform 1 0 78292 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_25_841
timestamp 1644511149
transform 1 0 78476 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_3
timestamp 1644511149
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_15
timestamp 1644511149
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1644511149
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_29
timestamp 1644511149
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_41
timestamp 1644511149
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_53
timestamp 1644511149
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_65
timestamp 1644511149
transform 1 0 7084 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_77
timestamp 1644511149
transform 1 0 8188 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1644511149
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_85
timestamp 1644511149
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_97
timestamp 1644511149
transform 1 0 10028 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_109
timestamp 1644511149
transform 1 0 11132 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_121
timestamp 1644511149
transform 1 0 12236 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_133
timestamp 1644511149
transform 1 0 13340 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_139
timestamp 1644511149
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_141
timestamp 1644511149
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_153
timestamp 1644511149
transform 1 0 15180 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_165
timestamp 1644511149
transform 1 0 16284 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_177
timestamp 1644511149
transform 1 0 17388 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_189
timestamp 1644511149
transform 1 0 18492 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_195
timestamp 1644511149
transform 1 0 19044 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_197
timestamp 1644511149
transform 1 0 19228 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_209
timestamp 1644511149
transform 1 0 20332 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_221
timestamp 1644511149
transform 1 0 21436 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_233
timestamp 1644511149
transform 1 0 22540 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_245
timestamp 1644511149
transform 1 0 23644 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_251
timestamp 1644511149
transform 1 0 24196 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_253
timestamp 1644511149
transform 1 0 24380 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_265
timestamp 1644511149
transform 1 0 25484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_277
timestamp 1644511149
transform 1 0 26588 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_289
timestamp 1644511149
transform 1 0 27692 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_301
timestamp 1644511149
transform 1 0 28796 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_307
timestamp 1644511149
transform 1 0 29348 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_309
timestamp 1644511149
transform 1 0 29532 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_321
timestamp 1644511149
transform 1 0 30636 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_333
timestamp 1644511149
transform 1 0 31740 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_345
timestamp 1644511149
transform 1 0 32844 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_357
timestamp 1644511149
transform 1 0 33948 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_363
timestamp 1644511149
transform 1 0 34500 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_365
timestamp 1644511149
transform 1 0 34684 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_377
timestamp 1644511149
transform 1 0 35788 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_389
timestamp 1644511149
transform 1 0 36892 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_401
timestamp 1644511149
transform 1 0 37996 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_413
timestamp 1644511149
transform 1 0 39100 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_419
timestamp 1644511149
transform 1 0 39652 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_421
timestamp 1644511149
transform 1 0 39836 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_433
timestamp 1644511149
transform 1 0 40940 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_445
timestamp 1644511149
transform 1 0 42044 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_457
timestamp 1644511149
transform 1 0 43148 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_469
timestamp 1644511149
transform 1 0 44252 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_475
timestamp 1644511149
transform 1 0 44804 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_477
timestamp 1644511149
transform 1 0 44988 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_489
timestamp 1644511149
transform 1 0 46092 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_501
timestamp 1644511149
transform 1 0 47196 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_513
timestamp 1644511149
transform 1 0 48300 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_525
timestamp 1644511149
transform 1 0 49404 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_531
timestamp 1644511149
transform 1 0 49956 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_533
timestamp 1644511149
transform 1 0 50140 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_545
timestamp 1644511149
transform 1 0 51244 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_557
timestamp 1644511149
transform 1 0 52348 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_569
timestamp 1644511149
transform 1 0 53452 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_581
timestamp 1644511149
transform 1 0 54556 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_587
timestamp 1644511149
transform 1 0 55108 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_589
timestamp 1644511149
transform 1 0 55292 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_601
timestamp 1644511149
transform 1 0 56396 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_613
timestamp 1644511149
transform 1 0 57500 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_625
timestamp 1644511149
transform 1 0 58604 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_637
timestamp 1644511149
transform 1 0 59708 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_643
timestamp 1644511149
transform 1 0 60260 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_645
timestamp 1644511149
transform 1 0 60444 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_657
timestamp 1644511149
transform 1 0 61548 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_669
timestamp 1644511149
transform 1 0 62652 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_681
timestamp 1644511149
transform 1 0 63756 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_693
timestamp 1644511149
transform 1 0 64860 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_699
timestamp 1644511149
transform 1 0 65412 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_701
timestamp 1644511149
transform 1 0 65596 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_713
timestamp 1644511149
transform 1 0 66700 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_725
timestamp 1644511149
transform 1 0 67804 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_737
timestamp 1644511149
transform 1 0 68908 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_749
timestamp 1644511149
transform 1 0 70012 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_755
timestamp 1644511149
transform 1 0 70564 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_757
timestamp 1644511149
transform 1 0 70748 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_769
timestamp 1644511149
transform 1 0 71852 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_781
timestamp 1644511149
transform 1 0 72956 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_793
timestamp 1644511149
transform 1 0 74060 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_805
timestamp 1644511149
transform 1 0 75164 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_811
timestamp 1644511149
transform 1 0 75716 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_813
timestamp 1644511149
transform 1 0 75900 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_825
timestamp 1644511149
transform 1 0 77004 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_833
timestamp 1644511149
transform 1 0 77740 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_838
timestamp 1644511149
transform 1 0 78200 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_27_3
timestamp 1644511149
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_15
timestamp 1644511149
transform 1 0 2484 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_27
timestamp 1644511149
transform 1 0 3588 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_39
timestamp 1644511149
transform 1 0 4692 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_51
timestamp 1644511149
transform 1 0 5796 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_55
timestamp 1644511149
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_57
timestamp 1644511149
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_69
timestamp 1644511149
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_81
timestamp 1644511149
transform 1 0 8556 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_93
timestamp 1644511149
transform 1 0 9660 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_105
timestamp 1644511149
transform 1 0 10764 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp 1644511149
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_113
timestamp 1644511149
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_125
timestamp 1644511149
transform 1 0 12604 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_137
timestamp 1644511149
transform 1 0 13708 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_149
timestamp 1644511149
transform 1 0 14812 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_161
timestamp 1644511149
transform 1 0 15916 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_167
timestamp 1644511149
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_169
timestamp 1644511149
transform 1 0 16652 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_181
timestamp 1644511149
transform 1 0 17756 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_193
timestamp 1644511149
transform 1 0 18860 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_205
timestamp 1644511149
transform 1 0 19964 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_217
timestamp 1644511149
transform 1 0 21068 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_223
timestamp 1644511149
transform 1 0 21620 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_225
timestamp 1644511149
transform 1 0 21804 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_237
timestamp 1644511149
transform 1 0 22908 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_249
timestamp 1644511149
transform 1 0 24012 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_261
timestamp 1644511149
transform 1 0 25116 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_273
timestamp 1644511149
transform 1 0 26220 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_279
timestamp 1644511149
transform 1 0 26772 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_281
timestamp 1644511149
transform 1 0 26956 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_293
timestamp 1644511149
transform 1 0 28060 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_305
timestamp 1644511149
transform 1 0 29164 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_317
timestamp 1644511149
transform 1 0 30268 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_329
timestamp 1644511149
transform 1 0 31372 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_335
timestamp 1644511149
transform 1 0 31924 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_337
timestamp 1644511149
transform 1 0 32108 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_349
timestamp 1644511149
transform 1 0 33212 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_361
timestamp 1644511149
transform 1 0 34316 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_373
timestamp 1644511149
transform 1 0 35420 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_385
timestamp 1644511149
transform 1 0 36524 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_391
timestamp 1644511149
transform 1 0 37076 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_393
timestamp 1644511149
transform 1 0 37260 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_405
timestamp 1644511149
transform 1 0 38364 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_417
timestamp 1644511149
transform 1 0 39468 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_429
timestamp 1644511149
transform 1 0 40572 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_441
timestamp 1644511149
transform 1 0 41676 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_447
timestamp 1644511149
transform 1 0 42228 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_449
timestamp 1644511149
transform 1 0 42412 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_461
timestamp 1644511149
transform 1 0 43516 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_473
timestamp 1644511149
transform 1 0 44620 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_485
timestamp 1644511149
transform 1 0 45724 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_497
timestamp 1644511149
transform 1 0 46828 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_503
timestamp 1644511149
transform 1 0 47380 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_505
timestamp 1644511149
transform 1 0 47564 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_517
timestamp 1644511149
transform 1 0 48668 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_529
timestamp 1644511149
transform 1 0 49772 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_541
timestamp 1644511149
transform 1 0 50876 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_553
timestamp 1644511149
transform 1 0 51980 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_559
timestamp 1644511149
transform 1 0 52532 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_561
timestamp 1644511149
transform 1 0 52716 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_573
timestamp 1644511149
transform 1 0 53820 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_585
timestamp 1644511149
transform 1 0 54924 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_597
timestamp 1644511149
transform 1 0 56028 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_609
timestamp 1644511149
transform 1 0 57132 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_615
timestamp 1644511149
transform 1 0 57684 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_617
timestamp 1644511149
transform 1 0 57868 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_629
timestamp 1644511149
transform 1 0 58972 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_641
timestamp 1644511149
transform 1 0 60076 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_653
timestamp 1644511149
transform 1 0 61180 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_665
timestamp 1644511149
transform 1 0 62284 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_671
timestamp 1644511149
transform 1 0 62836 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_673
timestamp 1644511149
transform 1 0 63020 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_685
timestamp 1644511149
transform 1 0 64124 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_697
timestamp 1644511149
transform 1 0 65228 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_709
timestamp 1644511149
transform 1 0 66332 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_721
timestamp 1644511149
transform 1 0 67436 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_727
timestamp 1644511149
transform 1 0 67988 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_729
timestamp 1644511149
transform 1 0 68172 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_741
timestamp 1644511149
transform 1 0 69276 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_753
timestamp 1644511149
transform 1 0 70380 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_765
timestamp 1644511149
transform 1 0 71484 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_777
timestamp 1644511149
transform 1 0 72588 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_783
timestamp 1644511149
transform 1 0 73140 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_785
timestamp 1644511149
transform 1 0 73324 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_797
timestamp 1644511149
transform 1 0 74428 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_809
timestamp 1644511149
transform 1 0 75532 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_821
timestamp 1644511149
transform 1 0 76636 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_833
timestamp 1644511149
transform 1 0 77740 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_839
timestamp 1644511149
transform 1 0 78292 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_841
timestamp 1644511149
transform 1 0 78476 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_3
timestamp 1644511149
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_15
timestamp 1644511149
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1644511149
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_29
timestamp 1644511149
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_41
timestamp 1644511149
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_53
timestamp 1644511149
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_65
timestamp 1644511149
transform 1 0 7084 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_77
timestamp 1644511149
transform 1 0 8188 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_83
timestamp 1644511149
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_85
timestamp 1644511149
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_97
timestamp 1644511149
transform 1 0 10028 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_109
timestamp 1644511149
transform 1 0 11132 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_121
timestamp 1644511149
transform 1 0 12236 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_133
timestamp 1644511149
transform 1 0 13340 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_139
timestamp 1644511149
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_141
timestamp 1644511149
transform 1 0 14076 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_153
timestamp 1644511149
transform 1 0 15180 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_165
timestamp 1644511149
transform 1 0 16284 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_177
timestamp 1644511149
transform 1 0 17388 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_189
timestamp 1644511149
transform 1 0 18492 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_195
timestamp 1644511149
transform 1 0 19044 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_197
timestamp 1644511149
transform 1 0 19228 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_209
timestamp 1644511149
transform 1 0 20332 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_221
timestamp 1644511149
transform 1 0 21436 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_233
timestamp 1644511149
transform 1 0 22540 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_245
timestamp 1644511149
transform 1 0 23644 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_251
timestamp 1644511149
transform 1 0 24196 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_253
timestamp 1644511149
transform 1 0 24380 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_265
timestamp 1644511149
transform 1 0 25484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_277
timestamp 1644511149
transform 1 0 26588 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_289
timestamp 1644511149
transform 1 0 27692 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_301
timestamp 1644511149
transform 1 0 28796 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_307
timestamp 1644511149
transform 1 0 29348 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_309
timestamp 1644511149
transform 1 0 29532 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_321
timestamp 1644511149
transform 1 0 30636 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_333
timestamp 1644511149
transform 1 0 31740 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_345
timestamp 1644511149
transform 1 0 32844 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_357
timestamp 1644511149
transform 1 0 33948 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_363
timestamp 1644511149
transform 1 0 34500 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_365
timestamp 1644511149
transform 1 0 34684 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_377
timestamp 1644511149
transform 1 0 35788 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_389
timestamp 1644511149
transform 1 0 36892 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_401
timestamp 1644511149
transform 1 0 37996 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_413
timestamp 1644511149
transform 1 0 39100 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_419
timestamp 1644511149
transform 1 0 39652 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_421
timestamp 1644511149
transform 1 0 39836 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_433
timestamp 1644511149
transform 1 0 40940 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_445
timestamp 1644511149
transform 1 0 42044 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_457
timestamp 1644511149
transform 1 0 43148 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_469
timestamp 1644511149
transform 1 0 44252 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_475
timestamp 1644511149
transform 1 0 44804 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_477
timestamp 1644511149
transform 1 0 44988 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_489
timestamp 1644511149
transform 1 0 46092 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_501
timestamp 1644511149
transform 1 0 47196 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_513
timestamp 1644511149
transform 1 0 48300 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_525
timestamp 1644511149
transform 1 0 49404 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_531
timestamp 1644511149
transform 1 0 49956 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_533
timestamp 1644511149
transform 1 0 50140 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_545
timestamp 1644511149
transform 1 0 51244 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_557
timestamp 1644511149
transform 1 0 52348 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_569
timestamp 1644511149
transform 1 0 53452 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_581
timestamp 1644511149
transform 1 0 54556 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_587
timestamp 1644511149
transform 1 0 55108 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_589
timestamp 1644511149
transform 1 0 55292 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_601
timestamp 1644511149
transform 1 0 56396 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_613
timestamp 1644511149
transform 1 0 57500 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_625
timestamp 1644511149
transform 1 0 58604 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_637
timestamp 1644511149
transform 1 0 59708 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_643
timestamp 1644511149
transform 1 0 60260 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_645
timestamp 1644511149
transform 1 0 60444 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_657
timestamp 1644511149
transform 1 0 61548 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_669
timestamp 1644511149
transform 1 0 62652 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_681
timestamp 1644511149
transform 1 0 63756 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_693
timestamp 1644511149
transform 1 0 64860 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_699
timestamp 1644511149
transform 1 0 65412 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_701
timestamp 1644511149
transform 1 0 65596 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_713
timestamp 1644511149
transform 1 0 66700 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_725
timestamp 1644511149
transform 1 0 67804 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_737
timestamp 1644511149
transform 1 0 68908 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_749
timestamp 1644511149
transform 1 0 70012 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_755
timestamp 1644511149
transform 1 0 70564 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_757
timestamp 1644511149
transform 1 0 70748 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_769
timestamp 1644511149
transform 1 0 71852 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_781
timestamp 1644511149
transform 1 0 72956 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_793
timestamp 1644511149
transform 1 0 74060 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_805
timestamp 1644511149
transform 1 0 75164 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_811
timestamp 1644511149
transform 1 0 75716 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_813
timestamp 1644511149
transform 1 0 75900 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_825
timestamp 1644511149
transform 1 0 77004 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_837
timestamp 1644511149
transform 1 0 78108 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_841
timestamp 1644511149
transform 1 0 78476 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_3
timestamp 1644511149
transform 1 0 1380 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_15
timestamp 1644511149
transform 1 0 2484 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_27
timestamp 1644511149
transform 1 0 3588 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_39
timestamp 1644511149
transform 1 0 4692 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_51
timestamp 1644511149
transform 1 0 5796 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_55
timestamp 1644511149
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_57
timestamp 1644511149
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_69
timestamp 1644511149
transform 1 0 7452 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_81
timestamp 1644511149
transform 1 0 8556 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_93
timestamp 1644511149
transform 1 0 9660 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_105
timestamp 1644511149
transform 1 0 10764 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_111
timestamp 1644511149
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_113
timestamp 1644511149
transform 1 0 11500 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_125
timestamp 1644511149
transform 1 0 12604 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_137
timestamp 1644511149
transform 1 0 13708 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_149
timestamp 1644511149
transform 1 0 14812 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_161
timestamp 1644511149
transform 1 0 15916 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_167
timestamp 1644511149
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_169
timestamp 1644511149
transform 1 0 16652 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_181
timestamp 1644511149
transform 1 0 17756 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_193
timestamp 1644511149
transform 1 0 18860 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_205
timestamp 1644511149
transform 1 0 19964 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_217
timestamp 1644511149
transform 1 0 21068 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_223
timestamp 1644511149
transform 1 0 21620 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_225
timestamp 1644511149
transform 1 0 21804 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_237
timestamp 1644511149
transform 1 0 22908 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_249
timestamp 1644511149
transform 1 0 24012 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_261
timestamp 1644511149
transform 1 0 25116 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_273
timestamp 1644511149
transform 1 0 26220 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_279
timestamp 1644511149
transform 1 0 26772 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_281
timestamp 1644511149
transform 1 0 26956 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_293
timestamp 1644511149
transform 1 0 28060 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_305
timestamp 1644511149
transform 1 0 29164 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_317
timestamp 1644511149
transform 1 0 30268 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_329
timestamp 1644511149
transform 1 0 31372 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_335
timestamp 1644511149
transform 1 0 31924 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_337
timestamp 1644511149
transform 1 0 32108 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_349
timestamp 1644511149
transform 1 0 33212 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_361
timestamp 1644511149
transform 1 0 34316 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_373
timestamp 1644511149
transform 1 0 35420 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_385
timestamp 1644511149
transform 1 0 36524 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_391
timestamp 1644511149
transform 1 0 37076 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_393
timestamp 1644511149
transform 1 0 37260 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_405
timestamp 1644511149
transform 1 0 38364 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_417
timestamp 1644511149
transform 1 0 39468 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_429
timestamp 1644511149
transform 1 0 40572 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_441
timestamp 1644511149
transform 1 0 41676 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_447
timestamp 1644511149
transform 1 0 42228 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_449
timestamp 1644511149
transform 1 0 42412 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_461
timestamp 1644511149
transform 1 0 43516 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_473
timestamp 1644511149
transform 1 0 44620 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_485
timestamp 1644511149
transform 1 0 45724 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_497
timestamp 1644511149
transform 1 0 46828 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_503
timestamp 1644511149
transform 1 0 47380 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_505
timestamp 1644511149
transform 1 0 47564 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_517
timestamp 1644511149
transform 1 0 48668 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_529
timestamp 1644511149
transform 1 0 49772 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_541
timestamp 1644511149
transform 1 0 50876 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_553
timestamp 1644511149
transform 1 0 51980 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_559
timestamp 1644511149
transform 1 0 52532 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_561
timestamp 1644511149
transform 1 0 52716 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_573
timestamp 1644511149
transform 1 0 53820 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_585
timestamp 1644511149
transform 1 0 54924 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_597
timestamp 1644511149
transform 1 0 56028 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_609
timestamp 1644511149
transform 1 0 57132 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_615
timestamp 1644511149
transform 1 0 57684 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_617
timestamp 1644511149
transform 1 0 57868 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_629
timestamp 1644511149
transform 1 0 58972 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_641
timestamp 1644511149
transform 1 0 60076 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_653
timestamp 1644511149
transform 1 0 61180 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_665
timestamp 1644511149
transform 1 0 62284 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_671
timestamp 1644511149
transform 1 0 62836 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_673
timestamp 1644511149
transform 1 0 63020 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_685
timestamp 1644511149
transform 1 0 64124 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_697
timestamp 1644511149
transform 1 0 65228 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_709
timestamp 1644511149
transform 1 0 66332 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_721
timestamp 1644511149
transform 1 0 67436 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_727
timestamp 1644511149
transform 1 0 67988 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_729
timestamp 1644511149
transform 1 0 68172 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_741
timestamp 1644511149
transform 1 0 69276 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_753
timestamp 1644511149
transform 1 0 70380 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_765
timestamp 1644511149
transform 1 0 71484 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_777
timestamp 1644511149
transform 1 0 72588 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_783
timestamp 1644511149
transform 1 0 73140 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_785
timestamp 1644511149
transform 1 0 73324 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_797
timestamp 1644511149
transform 1 0 74428 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_809
timestamp 1644511149
transform 1 0 75532 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_821
timestamp 1644511149
transform 1 0 76636 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_833
timestamp 1644511149
transform 1 0 77740 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_839
timestamp 1644511149
transform 1 0 78292 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_29_841
timestamp 1644511149
transform 1 0 78476 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_3
timestamp 1644511149
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_15
timestamp 1644511149
transform 1 0 2484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 1644511149
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_29
timestamp 1644511149
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_41
timestamp 1644511149
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_53
timestamp 1644511149
transform 1 0 5980 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_65
timestamp 1644511149
transform 1 0 7084 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_77
timestamp 1644511149
transform 1 0 8188 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp 1644511149
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_85
timestamp 1644511149
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_97
timestamp 1644511149
transform 1 0 10028 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_109
timestamp 1644511149
transform 1 0 11132 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_121
timestamp 1644511149
transform 1 0 12236 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_133
timestamp 1644511149
transform 1 0 13340 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_139
timestamp 1644511149
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_141
timestamp 1644511149
transform 1 0 14076 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_153
timestamp 1644511149
transform 1 0 15180 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_165
timestamp 1644511149
transform 1 0 16284 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_177
timestamp 1644511149
transform 1 0 17388 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_189
timestamp 1644511149
transform 1 0 18492 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_195
timestamp 1644511149
transform 1 0 19044 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_197
timestamp 1644511149
transform 1 0 19228 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_209
timestamp 1644511149
transform 1 0 20332 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_221
timestamp 1644511149
transform 1 0 21436 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_233
timestamp 1644511149
transform 1 0 22540 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_245
timestamp 1644511149
transform 1 0 23644 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_251
timestamp 1644511149
transform 1 0 24196 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_253
timestamp 1644511149
transform 1 0 24380 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_265
timestamp 1644511149
transform 1 0 25484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_277
timestamp 1644511149
transform 1 0 26588 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_289
timestamp 1644511149
transform 1 0 27692 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_301
timestamp 1644511149
transform 1 0 28796 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_307
timestamp 1644511149
transform 1 0 29348 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_309
timestamp 1644511149
transform 1 0 29532 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_321
timestamp 1644511149
transform 1 0 30636 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_333
timestamp 1644511149
transform 1 0 31740 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_345
timestamp 1644511149
transform 1 0 32844 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_357
timestamp 1644511149
transform 1 0 33948 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_363
timestamp 1644511149
transform 1 0 34500 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_365
timestamp 1644511149
transform 1 0 34684 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_377
timestamp 1644511149
transform 1 0 35788 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_389
timestamp 1644511149
transform 1 0 36892 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_401
timestamp 1644511149
transform 1 0 37996 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_413
timestamp 1644511149
transform 1 0 39100 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_419
timestamp 1644511149
transform 1 0 39652 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_421
timestamp 1644511149
transform 1 0 39836 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_433
timestamp 1644511149
transform 1 0 40940 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_445
timestamp 1644511149
transform 1 0 42044 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_457
timestamp 1644511149
transform 1 0 43148 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_469
timestamp 1644511149
transform 1 0 44252 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_475
timestamp 1644511149
transform 1 0 44804 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_477
timestamp 1644511149
transform 1 0 44988 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_489
timestamp 1644511149
transform 1 0 46092 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_501
timestamp 1644511149
transform 1 0 47196 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_513
timestamp 1644511149
transform 1 0 48300 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_525
timestamp 1644511149
transform 1 0 49404 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_531
timestamp 1644511149
transform 1 0 49956 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_533
timestamp 1644511149
transform 1 0 50140 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_545
timestamp 1644511149
transform 1 0 51244 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_557
timestamp 1644511149
transform 1 0 52348 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_569
timestamp 1644511149
transform 1 0 53452 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_581
timestamp 1644511149
transform 1 0 54556 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_587
timestamp 1644511149
transform 1 0 55108 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_589
timestamp 1644511149
transform 1 0 55292 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_601
timestamp 1644511149
transform 1 0 56396 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_613
timestamp 1644511149
transform 1 0 57500 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_625
timestamp 1644511149
transform 1 0 58604 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_637
timestamp 1644511149
transform 1 0 59708 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_643
timestamp 1644511149
transform 1 0 60260 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_645
timestamp 1644511149
transform 1 0 60444 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_657
timestamp 1644511149
transform 1 0 61548 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_669
timestamp 1644511149
transform 1 0 62652 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_681
timestamp 1644511149
transform 1 0 63756 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_693
timestamp 1644511149
transform 1 0 64860 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_699
timestamp 1644511149
transform 1 0 65412 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_701
timestamp 1644511149
transform 1 0 65596 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_713
timestamp 1644511149
transform 1 0 66700 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_725
timestamp 1644511149
transform 1 0 67804 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_737
timestamp 1644511149
transform 1 0 68908 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_749
timestamp 1644511149
transform 1 0 70012 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_755
timestamp 1644511149
transform 1 0 70564 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_757
timestamp 1644511149
transform 1 0 70748 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_769
timestamp 1644511149
transform 1 0 71852 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_781
timestamp 1644511149
transform 1 0 72956 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_793
timestamp 1644511149
transform 1 0 74060 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_805
timestamp 1644511149
transform 1 0 75164 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_811
timestamp 1644511149
transform 1 0 75716 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_813
timestamp 1644511149
transform 1 0 75900 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_825
timestamp 1644511149
transform 1 0 77004 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_837
timestamp 1644511149
transform 1 0 78108 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_841
timestamp 1644511149
transform 1 0 78476 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_7
timestamp 1644511149
transform 1 0 1748 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_19
timestamp 1644511149
transform 1 0 2852 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_31
timestamp 1644511149
transform 1 0 3956 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_43
timestamp 1644511149
transform 1 0 5060 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_31_55
timestamp 1644511149
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_57
timestamp 1644511149
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_69
timestamp 1644511149
transform 1 0 7452 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_81
timestamp 1644511149
transform 1 0 8556 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_93
timestamp 1644511149
transform 1 0 9660 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_105
timestamp 1644511149
transform 1 0 10764 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_111
timestamp 1644511149
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_113
timestamp 1644511149
transform 1 0 11500 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_125
timestamp 1644511149
transform 1 0 12604 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_137
timestamp 1644511149
transform 1 0 13708 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_149
timestamp 1644511149
transform 1 0 14812 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_161
timestamp 1644511149
transform 1 0 15916 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_167
timestamp 1644511149
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_169
timestamp 1644511149
transform 1 0 16652 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_181
timestamp 1644511149
transform 1 0 17756 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_193
timestamp 1644511149
transform 1 0 18860 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_205
timestamp 1644511149
transform 1 0 19964 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_217
timestamp 1644511149
transform 1 0 21068 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_223
timestamp 1644511149
transform 1 0 21620 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_225
timestamp 1644511149
transform 1 0 21804 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_237
timestamp 1644511149
transform 1 0 22908 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_249
timestamp 1644511149
transform 1 0 24012 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_261
timestamp 1644511149
transform 1 0 25116 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_273
timestamp 1644511149
transform 1 0 26220 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_279
timestamp 1644511149
transform 1 0 26772 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_281
timestamp 1644511149
transform 1 0 26956 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_293
timestamp 1644511149
transform 1 0 28060 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_305
timestamp 1644511149
transform 1 0 29164 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_317
timestamp 1644511149
transform 1 0 30268 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_329
timestamp 1644511149
transform 1 0 31372 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_335
timestamp 1644511149
transform 1 0 31924 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_337
timestamp 1644511149
transform 1 0 32108 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_349
timestamp 1644511149
transform 1 0 33212 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_361
timestamp 1644511149
transform 1 0 34316 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_373
timestamp 1644511149
transform 1 0 35420 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_385
timestamp 1644511149
transform 1 0 36524 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_391
timestamp 1644511149
transform 1 0 37076 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_393
timestamp 1644511149
transform 1 0 37260 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_405
timestamp 1644511149
transform 1 0 38364 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_417
timestamp 1644511149
transform 1 0 39468 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_429
timestamp 1644511149
transform 1 0 40572 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_441
timestamp 1644511149
transform 1 0 41676 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_447
timestamp 1644511149
transform 1 0 42228 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_449
timestamp 1644511149
transform 1 0 42412 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_461
timestamp 1644511149
transform 1 0 43516 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_473
timestamp 1644511149
transform 1 0 44620 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_485
timestamp 1644511149
transform 1 0 45724 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_497
timestamp 1644511149
transform 1 0 46828 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_503
timestamp 1644511149
transform 1 0 47380 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_505
timestamp 1644511149
transform 1 0 47564 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_517
timestamp 1644511149
transform 1 0 48668 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_529
timestamp 1644511149
transform 1 0 49772 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_541
timestamp 1644511149
transform 1 0 50876 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_553
timestamp 1644511149
transform 1 0 51980 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_559
timestamp 1644511149
transform 1 0 52532 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_561
timestamp 1644511149
transform 1 0 52716 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_573
timestamp 1644511149
transform 1 0 53820 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_585
timestamp 1644511149
transform 1 0 54924 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_597
timestamp 1644511149
transform 1 0 56028 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_609
timestamp 1644511149
transform 1 0 57132 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_615
timestamp 1644511149
transform 1 0 57684 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_617
timestamp 1644511149
transform 1 0 57868 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_629
timestamp 1644511149
transform 1 0 58972 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_641
timestamp 1644511149
transform 1 0 60076 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_653
timestamp 1644511149
transform 1 0 61180 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_665
timestamp 1644511149
transform 1 0 62284 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_671
timestamp 1644511149
transform 1 0 62836 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_673
timestamp 1644511149
transform 1 0 63020 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_685
timestamp 1644511149
transform 1 0 64124 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_697
timestamp 1644511149
transform 1 0 65228 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_709
timestamp 1644511149
transform 1 0 66332 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_721
timestamp 1644511149
transform 1 0 67436 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_727
timestamp 1644511149
transform 1 0 67988 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_729
timestamp 1644511149
transform 1 0 68172 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_741
timestamp 1644511149
transform 1 0 69276 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_753
timestamp 1644511149
transform 1 0 70380 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_765
timestamp 1644511149
transform 1 0 71484 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_777
timestamp 1644511149
transform 1 0 72588 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_783
timestamp 1644511149
transform 1 0 73140 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_785
timestamp 1644511149
transform 1 0 73324 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_797
timestamp 1644511149
transform 1 0 74428 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_809
timestamp 1644511149
transform 1 0 75532 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_821
timestamp 1644511149
transform 1 0 76636 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_833
timestamp 1644511149
transform 1 0 77740 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_839
timestamp 1644511149
transform 1 0 78292 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_31_841
timestamp 1644511149
transform 1 0 78476 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_3
timestamp 1644511149
transform 1 0 1380 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_15
timestamp 1644511149
transform 1 0 2484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1644511149
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_29
timestamp 1644511149
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_41
timestamp 1644511149
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_53
timestamp 1644511149
transform 1 0 5980 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_65
timestamp 1644511149
transform 1 0 7084 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_77
timestamp 1644511149
transform 1 0 8188 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_83
timestamp 1644511149
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_85
timestamp 1644511149
transform 1 0 8924 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_97
timestamp 1644511149
transform 1 0 10028 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_109
timestamp 1644511149
transform 1 0 11132 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_121
timestamp 1644511149
transform 1 0 12236 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_133
timestamp 1644511149
transform 1 0 13340 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_139
timestamp 1644511149
transform 1 0 13892 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_141
timestamp 1644511149
transform 1 0 14076 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_153
timestamp 1644511149
transform 1 0 15180 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_165
timestamp 1644511149
transform 1 0 16284 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_177
timestamp 1644511149
transform 1 0 17388 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_189
timestamp 1644511149
transform 1 0 18492 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_195
timestamp 1644511149
transform 1 0 19044 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_197
timestamp 1644511149
transform 1 0 19228 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_209
timestamp 1644511149
transform 1 0 20332 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_221
timestamp 1644511149
transform 1 0 21436 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_233
timestamp 1644511149
transform 1 0 22540 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_245
timestamp 1644511149
transform 1 0 23644 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_251
timestamp 1644511149
transform 1 0 24196 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_253
timestamp 1644511149
transform 1 0 24380 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_265
timestamp 1644511149
transform 1 0 25484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_277
timestamp 1644511149
transform 1 0 26588 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_289
timestamp 1644511149
transform 1 0 27692 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_301
timestamp 1644511149
transform 1 0 28796 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_307
timestamp 1644511149
transform 1 0 29348 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_309
timestamp 1644511149
transform 1 0 29532 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_321
timestamp 1644511149
transform 1 0 30636 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_333
timestamp 1644511149
transform 1 0 31740 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_345
timestamp 1644511149
transform 1 0 32844 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_357
timestamp 1644511149
transform 1 0 33948 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_363
timestamp 1644511149
transform 1 0 34500 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_365
timestamp 1644511149
transform 1 0 34684 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_377
timestamp 1644511149
transform 1 0 35788 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_389
timestamp 1644511149
transform 1 0 36892 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_401
timestamp 1644511149
transform 1 0 37996 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_413
timestamp 1644511149
transform 1 0 39100 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_419
timestamp 1644511149
transform 1 0 39652 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_421
timestamp 1644511149
transform 1 0 39836 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_433
timestamp 1644511149
transform 1 0 40940 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_445
timestamp 1644511149
transform 1 0 42044 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_457
timestamp 1644511149
transform 1 0 43148 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_469
timestamp 1644511149
transform 1 0 44252 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_475
timestamp 1644511149
transform 1 0 44804 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_477
timestamp 1644511149
transform 1 0 44988 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_489
timestamp 1644511149
transform 1 0 46092 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_501
timestamp 1644511149
transform 1 0 47196 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_513
timestamp 1644511149
transform 1 0 48300 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_525
timestamp 1644511149
transform 1 0 49404 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_531
timestamp 1644511149
transform 1 0 49956 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_533
timestamp 1644511149
transform 1 0 50140 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_545
timestamp 1644511149
transform 1 0 51244 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_557
timestamp 1644511149
transform 1 0 52348 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_569
timestamp 1644511149
transform 1 0 53452 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_581
timestamp 1644511149
transform 1 0 54556 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_587
timestamp 1644511149
transform 1 0 55108 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_589
timestamp 1644511149
transform 1 0 55292 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_601
timestamp 1644511149
transform 1 0 56396 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_613
timestamp 1644511149
transform 1 0 57500 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_625
timestamp 1644511149
transform 1 0 58604 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_637
timestamp 1644511149
transform 1 0 59708 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_643
timestamp 1644511149
transform 1 0 60260 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_645
timestamp 1644511149
transform 1 0 60444 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_657
timestamp 1644511149
transform 1 0 61548 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_669
timestamp 1644511149
transform 1 0 62652 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_681
timestamp 1644511149
transform 1 0 63756 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_693
timestamp 1644511149
transform 1 0 64860 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_699
timestamp 1644511149
transform 1 0 65412 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_701
timestamp 1644511149
transform 1 0 65596 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_713
timestamp 1644511149
transform 1 0 66700 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_725
timestamp 1644511149
transform 1 0 67804 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_737
timestamp 1644511149
transform 1 0 68908 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_749
timestamp 1644511149
transform 1 0 70012 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_755
timestamp 1644511149
transform 1 0 70564 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_757
timestamp 1644511149
transform 1 0 70748 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_769
timestamp 1644511149
transform 1 0 71852 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_781
timestamp 1644511149
transform 1 0 72956 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_793
timestamp 1644511149
transform 1 0 74060 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_805
timestamp 1644511149
transform 1 0 75164 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_811
timestamp 1644511149
transform 1 0 75716 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_813
timestamp 1644511149
transform 1 0 75900 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_825
timestamp 1644511149
transform 1 0 77004 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_837
timestamp 1644511149
transform 1 0 78108 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_841
timestamp 1644511149
transform 1 0 78476 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_3
timestamp 1644511149
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_15
timestamp 1644511149
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_27
timestamp 1644511149
transform 1 0 3588 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_39
timestamp 1644511149
transform 1 0 4692 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_51
timestamp 1644511149
transform 1 0 5796 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_55
timestamp 1644511149
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_57
timestamp 1644511149
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_69
timestamp 1644511149
transform 1 0 7452 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_81
timestamp 1644511149
transform 1 0 8556 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_93
timestamp 1644511149
transform 1 0 9660 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_105
timestamp 1644511149
transform 1 0 10764 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_111
timestamp 1644511149
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_113
timestamp 1644511149
transform 1 0 11500 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_125
timestamp 1644511149
transform 1 0 12604 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_137
timestamp 1644511149
transform 1 0 13708 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_149
timestamp 1644511149
transform 1 0 14812 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_161
timestamp 1644511149
transform 1 0 15916 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_167
timestamp 1644511149
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_169
timestamp 1644511149
transform 1 0 16652 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_181
timestamp 1644511149
transform 1 0 17756 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_193
timestamp 1644511149
transform 1 0 18860 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_205
timestamp 1644511149
transform 1 0 19964 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_217
timestamp 1644511149
transform 1 0 21068 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_223
timestamp 1644511149
transform 1 0 21620 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_225
timestamp 1644511149
transform 1 0 21804 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_237
timestamp 1644511149
transform 1 0 22908 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_249
timestamp 1644511149
transform 1 0 24012 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_261
timestamp 1644511149
transform 1 0 25116 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_273
timestamp 1644511149
transform 1 0 26220 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_279
timestamp 1644511149
transform 1 0 26772 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_281
timestamp 1644511149
transform 1 0 26956 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_293
timestamp 1644511149
transform 1 0 28060 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_305
timestamp 1644511149
transform 1 0 29164 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_317
timestamp 1644511149
transform 1 0 30268 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_329
timestamp 1644511149
transform 1 0 31372 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_335
timestamp 1644511149
transform 1 0 31924 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_337
timestamp 1644511149
transform 1 0 32108 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_349
timestamp 1644511149
transform 1 0 33212 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_361
timestamp 1644511149
transform 1 0 34316 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_373
timestamp 1644511149
transform 1 0 35420 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_385
timestamp 1644511149
transform 1 0 36524 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_391
timestamp 1644511149
transform 1 0 37076 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_393
timestamp 1644511149
transform 1 0 37260 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_405
timestamp 1644511149
transform 1 0 38364 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_417
timestamp 1644511149
transform 1 0 39468 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_429
timestamp 1644511149
transform 1 0 40572 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_441
timestamp 1644511149
transform 1 0 41676 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_447
timestamp 1644511149
transform 1 0 42228 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_449
timestamp 1644511149
transform 1 0 42412 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_461
timestamp 1644511149
transform 1 0 43516 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_473
timestamp 1644511149
transform 1 0 44620 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_485
timestamp 1644511149
transform 1 0 45724 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_497
timestamp 1644511149
transform 1 0 46828 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_503
timestamp 1644511149
transform 1 0 47380 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_505
timestamp 1644511149
transform 1 0 47564 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_517
timestamp 1644511149
transform 1 0 48668 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_529
timestamp 1644511149
transform 1 0 49772 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_541
timestamp 1644511149
transform 1 0 50876 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_553
timestamp 1644511149
transform 1 0 51980 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_559
timestamp 1644511149
transform 1 0 52532 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_561
timestamp 1644511149
transform 1 0 52716 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_573
timestamp 1644511149
transform 1 0 53820 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_585
timestamp 1644511149
transform 1 0 54924 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_597
timestamp 1644511149
transform 1 0 56028 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_609
timestamp 1644511149
transform 1 0 57132 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_615
timestamp 1644511149
transform 1 0 57684 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_617
timestamp 1644511149
transform 1 0 57868 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_629
timestamp 1644511149
transform 1 0 58972 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_641
timestamp 1644511149
transform 1 0 60076 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_653
timestamp 1644511149
transform 1 0 61180 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_665
timestamp 1644511149
transform 1 0 62284 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_671
timestamp 1644511149
transform 1 0 62836 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_673
timestamp 1644511149
transform 1 0 63020 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_685
timestamp 1644511149
transform 1 0 64124 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_697
timestamp 1644511149
transform 1 0 65228 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_709
timestamp 1644511149
transform 1 0 66332 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_721
timestamp 1644511149
transform 1 0 67436 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_727
timestamp 1644511149
transform 1 0 67988 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_729
timestamp 1644511149
transform 1 0 68172 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_741
timestamp 1644511149
transform 1 0 69276 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_753
timestamp 1644511149
transform 1 0 70380 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_765
timestamp 1644511149
transform 1 0 71484 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_777
timestamp 1644511149
transform 1 0 72588 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_783
timestamp 1644511149
transform 1 0 73140 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_785
timestamp 1644511149
transform 1 0 73324 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_797
timestamp 1644511149
transform 1 0 74428 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_809
timestamp 1644511149
transform 1 0 75532 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_821
timestamp 1644511149
transform 1 0 76636 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_833
timestamp 1644511149
transform 1 0 77740 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_839
timestamp 1644511149
transform 1 0 78292 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_33_841
timestamp 1644511149
transform 1 0 78476 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_3
timestamp 1644511149
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_15
timestamp 1644511149
transform 1 0 2484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1644511149
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_29
timestamp 1644511149
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_41
timestamp 1644511149
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_53
timestamp 1644511149
transform 1 0 5980 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_65
timestamp 1644511149
transform 1 0 7084 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_77
timestamp 1644511149
transform 1 0 8188 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_83
timestamp 1644511149
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_85
timestamp 1644511149
transform 1 0 8924 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_97
timestamp 1644511149
transform 1 0 10028 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_109
timestamp 1644511149
transform 1 0 11132 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_121
timestamp 1644511149
transform 1 0 12236 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_133
timestamp 1644511149
transform 1 0 13340 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_139
timestamp 1644511149
transform 1 0 13892 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_141
timestamp 1644511149
transform 1 0 14076 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_153
timestamp 1644511149
transform 1 0 15180 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_165
timestamp 1644511149
transform 1 0 16284 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_177
timestamp 1644511149
transform 1 0 17388 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_189
timestamp 1644511149
transform 1 0 18492 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_195
timestamp 1644511149
transform 1 0 19044 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_197
timestamp 1644511149
transform 1 0 19228 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_209
timestamp 1644511149
transform 1 0 20332 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_221
timestamp 1644511149
transform 1 0 21436 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_233
timestamp 1644511149
transform 1 0 22540 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_245
timestamp 1644511149
transform 1 0 23644 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_251
timestamp 1644511149
transform 1 0 24196 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_253
timestamp 1644511149
transform 1 0 24380 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_265
timestamp 1644511149
transform 1 0 25484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_277
timestamp 1644511149
transform 1 0 26588 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_289
timestamp 1644511149
transform 1 0 27692 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_301
timestamp 1644511149
transform 1 0 28796 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_307
timestamp 1644511149
transform 1 0 29348 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_309
timestamp 1644511149
transform 1 0 29532 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_321
timestamp 1644511149
transform 1 0 30636 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_333
timestamp 1644511149
transform 1 0 31740 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_345
timestamp 1644511149
transform 1 0 32844 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_357
timestamp 1644511149
transform 1 0 33948 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_363
timestamp 1644511149
transform 1 0 34500 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_365
timestamp 1644511149
transform 1 0 34684 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_377
timestamp 1644511149
transform 1 0 35788 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_389
timestamp 1644511149
transform 1 0 36892 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_401
timestamp 1644511149
transform 1 0 37996 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_413
timestamp 1644511149
transform 1 0 39100 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_419
timestamp 1644511149
transform 1 0 39652 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_421
timestamp 1644511149
transform 1 0 39836 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_433
timestamp 1644511149
transform 1 0 40940 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_445
timestamp 1644511149
transform 1 0 42044 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_457
timestamp 1644511149
transform 1 0 43148 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_469
timestamp 1644511149
transform 1 0 44252 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_475
timestamp 1644511149
transform 1 0 44804 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_477
timestamp 1644511149
transform 1 0 44988 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_489
timestamp 1644511149
transform 1 0 46092 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_501
timestamp 1644511149
transform 1 0 47196 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_513
timestamp 1644511149
transform 1 0 48300 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_525
timestamp 1644511149
transform 1 0 49404 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_531
timestamp 1644511149
transform 1 0 49956 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_533
timestamp 1644511149
transform 1 0 50140 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_545
timestamp 1644511149
transform 1 0 51244 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_557
timestamp 1644511149
transform 1 0 52348 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_569
timestamp 1644511149
transform 1 0 53452 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_581
timestamp 1644511149
transform 1 0 54556 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_587
timestamp 1644511149
transform 1 0 55108 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_589
timestamp 1644511149
transform 1 0 55292 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_601
timestamp 1644511149
transform 1 0 56396 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_613
timestamp 1644511149
transform 1 0 57500 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_625
timestamp 1644511149
transform 1 0 58604 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_637
timestamp 1644511149
transform 1 0 59708 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_643
timestamp 1644511149
transform 1 0 60260 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_645
timestamp 1644511149
transform 1 0 60444 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_657
timestamp 1644511149
transform 1 0 61548 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_669
timestamp 1644511149
transform 1 0 62652 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_681
timestamp 1644511149
transform 1 0 63756 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_693
timestamp 1644511149
transform 1 0 64860 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_699
timestamp 1644511149
transform 1 0 65412 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_701
timestamp 1644511149
transform 1 0 65596 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_713
timestamp 1644511149
transform 1 0 66700 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_725
timestamp 1644511149
transform 1 0 67804 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_737
timestamp 1644511149
transform 1 0 68908 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_749
timestamp 1644511149
transform 1 0 70012 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_755
timestamp 1644511149
transform 1 0 70564 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_757
timestamp 1644511149
transform 1 0 70748 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_769
timestamp 1644511149
transform 1 0 71852 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_781
timestamp 1644511149
transform 1 0 72956 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_793
timestamp 1644511149
transform 1 0 74060 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_805
timestamp 1644511149
transform 1 0 75164 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_811
timestamp 1644511149
transform 1 0 75716 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_813
timestamp 1644511149
transform 1 0 75900 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_825
timestamp 1644511149
transform 1 0 77004 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_833
timestamp 1644511149
transform 1 0 77740 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_838
timestamp 1644511149
transform 1 0 78200 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_35_3
timestamp 1644511149
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_15
timestamp 1644511149
transform 1 0 2484 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_27
timestamp 1644511149
transform 1 0 3588 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_39
timestamp 1644511149
transform 1 0 4692 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_51
timestamp 1644511149
transform 1 0 5796 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_55
timestamp 1644511149
transform 1 0 6164 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_57
timestamp 1644511149
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_69
timestamp 1644511149
transform 1 0 7452 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_81
timestamp 1644511149
transform 1 0 8556 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_93
timestamp 1644511149
transform 1 0 9660 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_105
timestamp 1644511149
transform 1 0 10764 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_111
timestamp 1644511149
transform 1 0 11316 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_113
timestamp 1644511149
transform 1 0 11500 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_125
timestamp 1644511149
transform 1 0 12604 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_137
timestamp 1644511149
transform 1 0 13708 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_149
timestamp 1644511149
transform 1 0 14812 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_161
timestamp 1644511149
transform 1 0 15916 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_167
timestamp 1644511149
transform 1 0 16468 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_169
timestamp 1644511149
transform 1 0 16652 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_181
timestamp 1644511149
transform 1 0 17756 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_193
timestamp 1644511149
transform 1 0 18860 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_205
timestamp 1644511149
transform 1 0 19964 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_217
timestamp 1644511149
transform 1 0 21068 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_223
timestamp 1644511149
transform 1 0 21620 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_225
timestamp 1644511149
transform 1 0 21804 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_237
timestamp 1644511149
transform 1 0 22908 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_249
timestamp 1644511149
transform 1 0 24012 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_261
timestamp 1644511149
transform 1 0 25116 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_273
timestamp 1644511149
transform 1 0 26220 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_279
timestamp 1644511149
transform 1 0 26772 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_281
timestamp 1644511149
transform 1 0 26956 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_293
timestamp 1644511149
transform 1 0 28060 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_305
timestamp 1644511149
transform 1 0 29164 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_317
timestamp 1644511149
transform 1 0 30268 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_329
timestamp 1644511149
transform 1 0 31372 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_335
timestamp 1644511149
transform 1 0 31924 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_337
timestamp 1644511149
transform 1 0 32108 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_349
timestamp 1644511149
transform 1 0 33212 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_361
timestamp 1644511149
transform 1 0 34316 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_373
timestamp 1644511149
transform 1 0 35420 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_385
timestamp 1644511149
transform 1 0 36524 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_391
timestamp 1644511149
transform 1 0 37076 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_393
timestamp 1644511149
transform 1 0 37260 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_405
timestamp 1644511149
transform 1 0 38364 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_417
timestamp 1644511149
transform 1 0 39468 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_429
timestamp 1644511149
transform 1 0 40572 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_441
timestamp 1644511149
transform 1 0 41676 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_447
timestamp 1644511149
transform 1 0 42228 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_449
timestamp 1644511149
transform 1 0 42412 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_461
timestamp 1644511149
transform 1 0 43516 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_473
timestamp 1644511149
transform 1 0 44620 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_485
timestamp 1644511149
transform 1 0 45724 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_497
timestamp 1644511149
transform 1 0 46828 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_503
timestamp 1644511149
transform 1 0 47380 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_505
timestamp 1644511149
transform 1 0 47564 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_517
timestamp 1644511149
transform 1 0 48668 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_529
timestamp 1644511149
transform 1 0 49772 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_541
timestamp 1644511149
transform 1 0 50876 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_553
timestamp 1644511149
transform 1 0 51980 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_559
timestamp 1644511149
transform 1 0 52532 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_561
timestamp 1644511149
transform 1 0 52716 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_573
timestamp 1644511149
transform 1 0 53820 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_585
timestamp 1644511149
transform 1 0 54924 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_597
timestamp 1644511149
transform 1 0 56028 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_609
timestamp 1644511149
transform 1 0 57132 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_615
timestamp 1644511149
transform 1 0 57684 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_617
timestamp 1644511149
transform 1 0 57868 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_629
timestamp 1644511149
transform 1 0 58972 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_641
timestamp 1644511149
transform 1 0 60076 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_653
timestamp 1644511149
transform 1 0 61180 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_665
timestamp 1644511149
transform 1 0 62284 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_671
timestamp 1644511149
transform 1 0 62836 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_673
timestamp 1644511149
transform 1 0 63020 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_685
timestamp 1644511149
transform 1 0 64124 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_697
timestamp 1644511149
transform 1 0 65228 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_709
timestamp 1644511149
transform 1 0 66332 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_721
timestamp 1644511149
transform 1 0 67436 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_727
timestamp 1644511149
transform 1 0 67988 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_729
timestamp 1644511149
transform 1 0 68172 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_741
timestamp 1644511149
transform 1 0 69276 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_753
timestamp 1644511149
transform 1 0 70380 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_765
timestamp 1644511149
transform 1 0 71484 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_777
timestamp 1644511149
transform 1 0 72588 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_783
timestamp 1644511149
transform 1 0 73140 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_785
timestamp 1644511149
transform 1 0 73324 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_797
timestamp 1644511149
transform 1 0 74428 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_809
timestamp 1644511149
transform 1 0 75532 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_821
timestamp 1644511149
transform 1 0 76636 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_833
timestamp 1644511149
transform 1 0 77740 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_839
timestamp 1644511149
transform 1 0 78292 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_35_841
timestamp 1644511149
transform 1 0 78476 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_3
timestamp 1644511149
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_15
timestamp 1644511149
transform 1 0 2484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 1644511149
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_29
timestamp 1644511149
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_41
timestamp 1644511149
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_53
timestamp 1644511149
transform 1 0 5980 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_65
timestamp 1644511149
transform 1 0 7084 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_77
timestamp 1644511149
transform 1 0 8188 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_83
timestamp 1644511149
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_85
timestamp 1644511149
transform 1 0 8924 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_97
timestamp 1644511149
transform 1 0 10028 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_109
timestamp 1644511149
transform 1 0 11132 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_121
timestamp 1644511149
transform 1 0 12236 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_133
timestamp 1644511149
transform 1 0 13340 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_139
timestamp 1644511149
transform 1 0 13892 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_141
timestamp 1644511149
transform 1 0 14076 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_153
timestamp 1644511149
transform 1 0 15180 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_165
timestamp 1644511149
transform 1 0 16284 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_177
timestamp 1644511149
transform 1 0 17388 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_189
timestamp 1644511149
transform 1 0 18492 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_195
timestamp 1644511149
transform 1 0 19044 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_197
timestamp 1644511149
transform 1 0 19228 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_209
timestamp 1644511149
transform 1 0 20332 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_221
timestamp 1644511149
transform 1 0 21436 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_233
timestamp 1644511149
transform 1 0 22540 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_245
timestamp 1644511149
transform 1 0 23644 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_251
timestamp 1644511149
transform 1 0 24196 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_253
timestamp 1644511149
transform 1 0 24380 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_265
timestamp 1644511149
transform 1 0 25484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_277
timestamp 1644511149
transform 1 0 26588 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_289
timestamp 1644511149
transform 1 0 27692 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_301
timestamp 1644511149
transform 1 0 28796 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_307
timestamp 1644511149
transform 1 0 29348 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_309
timestamp 1644511149
transform 1 0 29532 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_321
timestamp 1644511149
transform 1 0 30636 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_333
timestamp 1644511149
transform 1 0 31740 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_345
timestamp 1644511149
transform 1 0 32844 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_357
timestamp 1644511149
transform 1 0 33948 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_363
timestamp 1644511149
transform 1 0 34500 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_365
timestamp 1644511149
transform 1 0 34684 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_377
timestamp 1644511149
transform 1 0 35788 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_389
timestamp 1644511149
transform 1 0 36892 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_401
timestamp 1644511149
transform 1 0 37996 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_413
timestamp 1644511149
transform 1 0 39100 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_419
timestamp 1644511149
transform 1 0 39652 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_421
timestamp 1644511149
transform 1 0 39836 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_433
timestamp 1644511149
transform 1 0 40940 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_445
timestamp 1644511149
transform 1 0 42044 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_457
timestamp 1644511149
transform 1 0 43148 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_469
timestamp 1644511149
transform 1 0 44252 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_475
timestamp 1644511149
transform 1 0 44804 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_477
timestamp 1644511149
transform 1 0 44988 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_489
timestamp 1644511149
transform 1 0 46092 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_501
timestamp 1644511149
transform 1 0 47196 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_513
timestamp 1644511149
transform 1 0 48300 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_525
timestamp 1644511149
transform 1 0 49404 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_531
timestamp 1644511149
transform 1 0 49956 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_533
timestamp 1644511149
transform 1 0 50140 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_545
timestamp 1644511149
transform 1 0 51244 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_557
timestamp 1644511149
transform 1 0 52348 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_569
timestamp 1644511149
transform 1 0 53452 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_581
timestamp 1644511149
transform 1 0 54556 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_587
timestamp 1644511149
transform 1 0 55108 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_589
timestamp 1644511149
transform 1 0 55292 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_601
timestamp 1644511149
transform 1 0 56396 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_613
timestamp 1644511149
transform 1 0 57500 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_625
timestamp 1644511149
transform 1 0 58604 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_637
timestamp 1644511149
transform 1 0 59708 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_643
timestamp 1644511149
transform 1 0 60260 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_645
timestamp 1644511149
transform 1 0 60444 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_657
timestamp 1644511149
transform 1 0 61548 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_669
timestamp 1644511149
transform 1 0 62652 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_681
timestamp 1644511149
transform 1 0 63756 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_693
timestamp 1644511149
transform 1 0 64860 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_699
timestamp 1644511149
transform 1 0 65412 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_701
timestamp 1644511149
transform 1 0 65596 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_713
timestamp 1644511149
transform 1 0 66700 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_725
timestamp 1644511149
transform 1 0 67804 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_737
timestamp 1644511149
transform 1 0 68908 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_749
timestamp 1644511149
transform 1 0 70012 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_755
timestamp 1644511149
transform 1 0 70564 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_757
timestamp 1644511149
transform 1 0 70748 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_769
timestamp 1644511149
transform 1 0 71852 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_781
timestamp 1644511149
transform 1 0 72956 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_793
timestamp 1644511149
transform 1 0 74060 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_805
timestamp 1644511149
transform 1 0 75164 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_811
timestamp 1644511149
transform 1 0 75716 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_813
timestamp 1644511149
transform 1 0 75900 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_825
timestamp 1644511149
transform 1 0 77004 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_837
timestamp 1644511149
transform 1 0 78108 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_841
timestamp 1644511149
transform 1 0 78476 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_3
timestamp 1644511149
transform 1 0 1380 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_15
timestamp 1644511149
transform 1 0 2484 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_27
timestamp 1644511149
transform 1 0 3588 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_39
timestamp 1644511149
transform 1 0 4692 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_51
timestamp 1644511149
transform 1 0 5796 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_55
timestamp 1644511149
transform 1 0 6164 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_57
timestamp 1644511149
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_69
timestamp 1644511149
transform 1 0 7452 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_81
timestamp 1644511149
transform 1 0 8556 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_93
timestamp 1644511149
transform 1 0 9660 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_105
timestamp 1644511149
transform 1 0 10764 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_111
timestamp 1644511149
transform 1 0 11316 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_113
timestamp 1644511149
transform 1 0 11500 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_125
timestamp 1644511149
transform 1 0 12604 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_137
timestamp 1644511149
transform 1 0 13708 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_149
timestamp 1644511149
transform 1 0 14812 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_161
timestamp 1644511149
transform 1 0 15916 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_167
timestamp 1644511149
transform 1 0 16468 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_169
timestamp 1644511149
transform 1 0 16652 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_181
timestamp 1644511149
transform 1 0 17756 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_193
timestamp 1644511149
transform 1 0 18860 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_205
timestamp 1644511149
transform 1 0 19964 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_217
timestamp 1644511149
transform 1 0 21068 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_223
timestamp 1644511149
transform 1 0 21620 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_225
timestamp 1644511149
transform 1 0 21804 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_237
timestamp 1644511149
transform 1 0 22908 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_249
timestamp 1644511149
transform 1 0 24012 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_261
timestamp 1644511149
transform 1 0 25116 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_273
timestamp 1644511149
transform 1 0 26220 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_279
timestamp 1644511149
transform 1 0 26772 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_281
timestamp 1644511149
transform 1 0 26956 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_293
timestamp 1644511149
transform 1 0 28060 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_305
timestamp 1644511149
transform 1 0 29164 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_317
timestamp 1644511149
transform 1 0 30268 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_329
timestamp 1644511149
transform 1 0 31372 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_335
timestamp 1644511149
transform 1 0 31924 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_337
timestamp 1644511149
transform 1 0 32108 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_349
timestamp 1644511149
transform 1 0 33212 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_361
timestamp 1644511149
transform 1 0 34316 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_373
timestamp 1644511149
transform 1 0 35420 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_385
timestamp 1644511149
transform 1 0 36524 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_391
timestamp 1644511149
transform 1 0 37076 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_393
timestamp 1644511149
transform 1 0 37260 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_405
timestamp 1644511149
transform 1 0 38364 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_417
timestamp 1644511149
transform 1 0 39468 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_429
timestamp 1644511149
transform 1 0 40572 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_441
timestamp 1644511149
transform 1 0 41676 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_447
timestamp 1644511149
transform 1 0 42228 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_449
timestamp 1644511149
transform 1 0 42412 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_461
timestamp 1644511149
transform 1 0 43516 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_473
timestamp 1644511149
transform 1 0 44620 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_485
timestamp 1644511149
transform 1 0 45724 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_497
timestamp 1644511149
transform 1 0 46828 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_503
timestamp 1644511149
transform 1 0 47380 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_505
timestamp 1644511149
transform 1 0 47564 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_517
timestamp 1644511149
transform 1 0 48668 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_529
timestamp 1644511149
transform 1 0 49772 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_541
timestamp 1644511149
transform 1 0 50876 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_553
timestamp 1644511149
transform 1 0 51980 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_559
timestamp 1644511149
transform 1 0 52532 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_561
timestamp 1644511149
transform 1 0 52716 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_573
timestamp 1644511149
transform 1 0 53820 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_585
timestamp 1644511149
transform 1 0 54924 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_597
timestamp 1644511149
transform 1 0 56028 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_609
timestamp 1644511149
transform 1 0 57132 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_615
timestamp 1644511149
transform 1 0 57684 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_617
timestamp 1644511149
transform 1 0 57868 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_629
timestamp 1644511149
transform 1 0 58972 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_641
timestamp 1644511149
transform 1 0 60076 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_653
timestamp 1644511149
transform 1 0 61180 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_665
timestamp 1644511149
transform 1 0 62284 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_671
timestamp 1644511149
transform 1 0 62836 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_673
timestamp 1644511149
transform 1 0 63020 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_685
timestamp 1644511149
transform 1 0 64124 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_697
timestamp 1644511149
transform 1 0 65228 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_709
timestamp 1644511149
transform 1 0 66332 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_721
timestamp 1644511149
transform 1 0 67436 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_727
timestamp 1644511149
transform 1 0 67988 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_729
timestamp 1644511149
transform 1 0 68172 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_741
timestamp 1644511149
transform 1 0 69276 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_753
timestamp 1644511149
transform 1 0 70380 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_765
timestamp 1644511149
transform 1 0 71484 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_777
timestamp 1644511149
transform 1 0 72588 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_783
timestamp 1644511149
transform 1 0 73140 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_785
timestamp 1644511149
transform 1 0 73324 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_797
timestamp 1644511149
transform 1 0 74428 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_809
timestamp 1644511149
transform 1 0 75532 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_821
timestamp 1644511149
transform 1 0 76636 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_833
timestamp 1644511149
transform 1 0 77740 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_839
timestamp 1644511149
transform 1 0 78292 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_37_841
timestamp 1644511149
transform 1 0 78476 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_3
timestamp 1644511149
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_15
timestamp 1644511149
transform 1 0 2484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 1644511149
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_29
timestamp 1644511149
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_41
timestamp 1644511149
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_53
timestamp 1644511149
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_65
timestamp 1644511149
transform 1 0 7084 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_77
timestamp 1644511149
transform 1 0 8188 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_83
timestamp 1644511149
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_85
timestamp 1644511149
transform 1 0 8924 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_97
timestamp 1644511149
transform 1 0 10028 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_109
timestamp 1644511149
transform 1 0 11132 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_121
timestamp 1644511149
transform 1 0 12236 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_133
timestamp 1644511149
transform 1 0 13340 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_139
timestamp 1644511149
transform 1 0 13892 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_141
timestamp 1644511149
transform 1 0 14076 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_153
timestamp 1644511149
transform 1 0 15180 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_165
timestamp 1644511149
transform 1 0 16284 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_177
timestamp 1644511149
transform 1 0 17388 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_189
timestamp 1644511149
transform 1 0 18492 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_195
timestamp 1644511149
transform 1 0 19044 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_197
timestamp 1644511149
transform 1 0 19228 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_209
timestamp 1644511149
transform 1 0 20332 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_221
timestamp 1644511149
transform 1 0 21436 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_233
timestamp 1644511149
transform 1 0 22540 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_245
timestamp 1644511149
transform 1 0 23644 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_251
timestamp 1644511149
transform 1 0 24196 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_253
timestamp 1644511149
transform 1 0 24380 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_265
timestamp 1644511149
transform 1 0 25484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_277
timestamp 1644511149
transform 1 0 26588 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_289
timestamp 1644511149
transform 1 0 27692 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_301
timestamp 1644511149
transform 1 0 28796 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_307
timestamp 1644511149
transform 1 0 29348 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_309
timestamp 1644511149
transform 1 0 29532 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_321
timestamp 1644511149
transform 1 0 30636 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_333
timestamp 1644511149
transform 1 0 31740 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_345
timestamp 1644511149
transform 1 0 32844 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_357
timestamp 1644511149
transform 1 0 33948 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_363
timestamp 1644511149
transform 1 0 34500 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_365
timestamp 1644511149
transform 1 0 34684 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_377
timestamp 1644511149
transform 1 0 35788 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_389
timestamp 1644511149
transform 1 0 36892 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_401
timestamp 1644511149
transform 1 0 37996 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_413
timestamp 1644511149
transform 1 0 39100 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_419
timestamp 1644511149
transform 1 0 39652 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_421
timestamp 1644511149
transform 1 0 39836 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_433
timestamp 1644511149
transform 1 0 40940 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_445
timestamp 1644511149
transform 1 0 42044 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_457
timestamp 1644511149
transform 1 0 43148 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_469
timestamp 1644511149
transform 1 0 44252 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_475
timestamp 1644511149
transform 1 0 44804 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_477
timestamp 1644511149
transform 1 0 44988 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_489
timestamp 1644511149
transform 1 0 46092 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_501
timestamp 1644511149
transform 1 0 47196 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_513
timestamp 1644511149
transform 1 0 48300 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_525
timestamp 1644511149
transform 1 0 49404 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_531
timestamp 1644511149
transform 1 0 49956 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_533
timestamp 1644511149
transform 1 0 50140 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_545
timestamp 1644511149
transform 1 0 51244 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_557
timestamp 1644511149
transform 1 0 52348 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_569
timestamp 1644511149
transform 1 0 53452 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_581
timestamp 1644511149
transform 1 0 54556 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_587
timestamp 1644511149
transform 1 0 55108 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_589
timestamp 1644511149
transform 1 0 55292 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_601
timestamp 1644511149
transform 1 0 56396 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_613
timestamp 1644511149
transform 1 0 57500 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_625
timestamp 1644511149
transform 1 0 58604 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_637
timestamp 1644511149
transform 1 0 59708 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_643
timestamp 1644511149
transform 1 0 60260 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_645
timestamp 1644511149
transform 1 0 60444 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_657
timestamp 1644511149
transform 1 0 61548 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_669
timestamp 1644511149
transform 1 0 62652 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_681
timestamp 1644511149
transform 1 0 63756 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_693
timestamp 1644511149
transform 1 0 64860 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_699
timestamp 1644511149
transform 1 0 65412 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_701
timestamp 1644511149
transform 1 0 65596 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_713
timestamp 1644511149
transform 1 0 66700 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_725
timestamp 1644511149
transform 1 0 67804 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_737
timestamp 1644511149
transform 1 0 68908 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_749
timestamp 1644511149
transform 1 0 70012 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_755
timestamp 1644511149
transform 1 0 70564 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_757
timestamp 1644511149
transform 1 0 70748 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_769
timestamp 1644511149
transform 1 0 71852 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_781
timestamp 1644511149
transform 1 0 72956 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_793
timestamp 1644511149
transform 1 0 74060 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_805
timestamp 1644511149
transform 1 0 75164 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_811
timestamp 1644511149
transform 1 0 75716 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_813
timestamp 1644511149
transform 1 0 75900 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_825
timestamp 1644511149
transform 1 0 77004 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_837
timestamp 1644511149
transform 1 0 78108 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_841
timestamp 1644511149
transform 1 0 78476 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_9
timestamp 1644511149
transform 1 0 1932 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_21
timestamp 1644511149
transform 1 0 3036 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_33
timestamp 1644511149
transform 1 0 4140 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_45
timestamp 1644511149
transform 1 0 5244 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_39_53
timestamp 1644511149
transform 1 0 5980 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_39_57
timestamp 1644511149
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_69
timestamp 1644511149
transform 1 0 7452 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_81
timestamp 1644511149
transform 1 0 8556 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_93
timestamp 1644511149
transform 1 0 9660 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_105
timestamp 1644511149
transform 1 0 10764 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_111
timestamp 1644511149
transform 1 0 11316 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_113
timestamp 1644511149
transform 1 0 11500 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_125
timestamp 1644511149
transform 1 0 12604 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_137
timestamp 1644511149
transform 1 0 13708 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_149
timestamp 1644511149
transform 1 0 14812 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_161
timestamp 1644511149
transform 1 0 15916 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_167
timestamp 1644511149
transform 1 0 16468 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_169
timestamp 1644511149
transform 1 0 16652 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_181
timestamp 1644511149
transform 1 0 17756 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_193
timestamp 1644511149
transform 1 0 18860 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_205
timestamp 1644511149
transform 1 0 19964 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_217
timestamp 1644511149
transform 1 0 21068 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_223
timestamp 1644511149
transform 1 0 21620 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_225
timestamp 1644511149
transform 1 0 21804 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_237
timestamp 1644511149
transform 1 0 22908 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_249
timestamp 1644511149
transform 1 0 24012 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_261
timestamp 1644511149
transform 1 0 25116 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_273
timestamp 1644511149
transform 1 0 26220 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_279
timestamp 1644511149
transform 1 0 26772 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_281
timestamp 1644511149
transform 1 0 26956 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_293
timestamp 1644511149
transform 1 0 28060 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_305
timestamp 1644511149
transform 1 0 29164 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_317
timestamp 1644511149
transform 1 0 30268 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_329
timestamp 1644511149
transform 1 0 31372 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_335
timestamp 1644511149
transform 1 0 31924 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_337
timestamp 1644511149
transform 1 0 32108 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_349
timestamp 1644511149
transform 1 0 33212 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_361
timestamp 1644511149
transform 1 0 34316 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_373
timestamp 1644511149
transform 1 0 35420 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_385
timestamp 1644511149
transform 1 0 36524 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_391
timestamp 1644511149
transform 1 0 37076 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_393
timestamp 1644511149
transform 1 0 37260 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_405
timestamp 1644511149
transform 1 0 38364 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_417
timestamp 1644511149
transform 1 0 39468 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_429
timestamp 1644511149
transform 1 0 40572 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_441
timestamp 1644511149
transform 1 0 41676 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_447
timestamp 1644511149
transform 1 0 42228 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_449
timestamp 1644511149
transform 1 0 42412 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_461
timestamp 1644511149
transform 1 0 43516 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_473
timestamp 1644511149
transform 1 0 44620 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_485
timestamp 1644511149
transform 1 0 45724 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_497
timestamp 1644511149
transform 1 0 46828 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_503
timestamp 1644511149
transform 1 0 47380 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_505
timestamp 1644511149
transform 1 0 47564 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_517
timestamp 1644511149
transform 1 0 48668 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_529
timestamp 1644511149
transform 1 0 49772 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_541
timestamp 1644511149
transform 1 0 50876 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_553
timestamp 1644511149
transform 1 0 51980 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_559
timestamp 1644511149
transform 1 0 52532 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_561
timestamp 1644511149
transform 1 0 52716 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_573
timestamp 1644511149
transform 1 0 53820 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_585
timestamp 1644511149
transform 1 0 54924 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_597
timestamp 1644511149
transform 1 0 56028 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_609
timestamp 1644511149
transform 1 0 57132 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_615
timestamp 1644511149
transform 1 0 57684 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_617
timestamp 1644511149
transform 1 0 57868 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_629
timestamp 1644511149
transform 1 0 58972 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_641
timestamp 1644511149
transform 1 0 60076 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_653
timestamp 1644511149
transform 1 0 61180 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_665
timestamp 1644511149
transform 1 0 62284 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_671
timestamp 1644511149
transform 1 0 62836 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_673
timestamp 1644511149
transform 1 0 63020 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_685
timestamp 1644511149
transform 1 0 64124 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_697
timestamp 1644511149
transform 1 0 65228 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_709
timestamp 1644511149
transform 1 0 66332 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_721
timestamp 1644511149
transform 1 0 67436 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_727
timestamp 1644511149
transform 1 0 67988 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_729
timestamp 1644511149
transform 1 0 68172 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_741
timestamp 1644511149
transform 1 0 69276 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_753
timestamp 1644511149
transform 1 0 70380 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_765
timestamp 1644511149
transform 1 0 71484 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_777
timestamp 1644511149
transform 1 0 72588 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_783
timestamp 1644511149
transform 1 0 73140 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_785
timestamp 1644511149
transform 1 0 73324 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_797
timestamp 1644511149
transform 1 0 74428 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_809
timestamp 1644511149
transform 1 0 75532 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_821
timestamp 1644511149
transform 1 0 76636 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_833
timestamp 1644511149
transform 1 0 77740 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_839
timestamp 1644511149
transform 1 0 78292 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_39_841
timestamp 1644511149
transform 1 0 78476 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_3
timestamp 1644511149
transform 1 0 1380 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_15
timestamp 1644511149
transform 1 0 2484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_27
timestamp 1644511149
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_29
timestamp 1644511149
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_41
timestamp 1644511149
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_53
timestamp 1644511149
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_65
timestamp 1644511149
transform 1 0 7084 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_77
timestamp 1644511149
transform 1 0 8188 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_83
timestamp 1644511149
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_85
timestamp 1644511149
transform 1 0 8924 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_97
timestamp 1644511149
transform 1 0 10028 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_109
timestamp 1644511149
transform 1 0 11132 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_121
timestamp 1644511149
transform 1 0 12236 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_133
timestamp 1644511149
transform 1 0 13340 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_139
timestamp 1644511149
transform 1 0 13892 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_141
timestamp 1644511149
transform 1 0 14076 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_153
timestamp 1644511149
transform 1 0 15180 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_165
timestamp 1644511149
transform 1 0 16284 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_177
timestamp 1644511149
transform 1 0 17388 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_189
timestamp 1644511149
transform 1 0 18492 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_195
timestamp 1644511149
transform 1 0 19044 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_197
timestamp 1644511149
transform 1 0 19228 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_209
timestamp 1644511149
transform 1 0 20332 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_221
timestamp 1644511149
transform 1 0 21436 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_233
timestamp 1644511149
transform 1 0 22540 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_245
timestamp 1644511149
transform 1 0 23644 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_251
timestamp 1644511149
transform 1 0 24196 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_253
timestamp 1644511149
transform 1 0 24380 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_265
timestamp 1644511149
transform 1 0 25484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_277
timestamp 1644511149
transform 1 0 26588 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_289
timestamp 1644511149
transform 1 0 27692 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_301
timestamp 1644511149
transform 1 0 28796 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_307
timestamp 1644511149
transform 1 0 29348 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_309
timestamp 1644511149
transform 1 0 29532 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_321
timestamp 1644511149
transform 1 0 30636 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_333
timestamp 1644511149
transform 1 0 31740 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_345
timestamp 1644511149
transform 1 0 32844 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_357
timestamp 1644511149
transform 1 0 33948 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_363
timestamp 1644511149
transform 1 0 34500 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_365
timestamp 1644511149
transform 1 0 34684 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_377
timestamp 1644511149
transform 1 0 35788 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_389
timestamp 1644511149
transform 1 0 36892 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_401
timestamp 1644511149
transform 1 0 37996 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_413
timestamp 1644511149
transform 1 0 39100 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_419
timestamp 1644511149
transform 1 0 39652 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_421
timestamp 1644511149
transform 1 0 39836 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_433
timestamp 1644511149
transform 1 0 40940 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_445
timestamp 1644511149
transform 1 0 42044 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_457
timestamp 1644511149
transform 1 0 43148 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_469
timestamp 1644511149
transform 1 0 44252 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_475
timestamp 1644511149
transform 1 0 44804 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_477
timestamp 1644511149
transform 1 0 44988 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_489
timestamp 1644511149
transform 1 0 46092 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_501
timestamp 1644511149
transform 1 0 47196 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_513
timestamp 1644511149
transform 1 0 48300 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_525
timestamp 1644511149
transform 1 0 49404 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_531
timestamp 1644511149
transform 1 0 49956 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_533
timestamp 1644511149
transform 1 0 50140 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_545
timestamp 1644511149
transform 1 0 51244 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_557
timestamp 1644511149
transform 1 0 52348 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_569
timestamp 1644511149
transform 1 0 53452 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_581
timestamp 1644511149
transform 1 0 54556 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_587
timestamp 1644511149
transform 1 0 55108 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_589
timestamp 1644511149
transform 1 0 55292 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_601
timestamp 1644511149
transform 1 0 56396 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_613
timestamp 1644511149
transform 1 0 57500 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_625
timestamp 1644511149
transform 1 0 58604 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_637
timestamp 1644511149
transform 1 0 59708 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_643
timestamp 1644511149
transform 1 0 60260 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_645
timestamp 1644511149
transform 1 0 60444 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_657
timestamp 1644511149
transform 1 0 61548 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_669
timestamp 1644511149
transform 1 0 62652 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_681
timestamp 1644511149
transform 1 0 63756 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_693
timestamp 1644511149
transform 1 0 64860 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_699
timestamp 1644511149
transform 1 0 65412 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_701
timestamp 1644511149
transform 1 0 65596 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_713
timestamp 1644511149
transform 1 0 66700 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_725
timestamp 1644511149
transform 1 0 67804 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_737
timestamp 1644511149
transform 1 0 68908 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_749
timestamp 1644511149
transform 1 0 70012 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_755
timestamp 1644511149
transform 1 0 70564 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_757
timestamp 1644511149
transform 1 0 70748 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_769
timestamp 1644511149
transform 1 0 71852 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_781
timestamp 1644511149
transform 1 0 72956 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_793
timestamp 1644511149
transform 1 0 74060 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_805
timestamp 1644511149
transform 1 0 75164 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_811
timestamp 1644511149
transform 1 0 75716 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_813
timestamp 1644511149
transform 1 0 75900 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_825
timestamp 1644511149
transform 1 0 77004 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_837
timestamp 1644511149
transform 1 0 78108 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_841
timestamp 1644511149
transform 1 0 78476 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_3
timestamp 1644511149
transform 1 0 1380 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_15
timestamp 1644511149
transform 1 0 2484 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_27
timestamp 1644511149
transform 1 0 3588 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_39
timestamp 1644511149
transform 1 0 4692 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_51
timestamp 1644511149
transform 1 0 5796 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_55
timestamp 1644511149
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_57
timestamp 1644511149
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_69
timestamp 1644511149
transform 1 0 7452 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_81
timestamp 1644511149
transform 1 0 8556 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_93
timestamp 1644511149
transform 1 0 9660 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_105
timestamp 1644511149
transform 1 0 10764 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_111
timestamp 1644511149
transform 1 0 11316 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_113
timestamp 1644511149
transform 1 0 11500 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_125
timestamp 1644511149
transform 1 0 12604 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_137
timestamp 1644511149
transform 1 0 13708 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_149
timestamp 1644511149
transform 1 0 14812 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_161
timestamp 1644511149
transform 1 0 15916 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_167
timestamp 1644511149
transform 1 0 16468 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_169
timestamp 1644511149
transform 1 0 16652 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_181
timestamp 1644511149
transform 1 0 17756 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_193
timestamp 1644511149
transform 1 0 18860 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_205
timestamp 1644511149
transform 1 0 19964 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_217
timestamp 1644511149
transform 1 0 21068 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_223
timestamp 1644511149
transform 1 0 21620 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_225
timestamp 1644511149
transform 1 0 21804 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_237
timestamp 1644511149
transform 1 0 22908 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_249
timestamp 1644511149
transform 1 0 24012 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_261
timestamp 1644511149
transform 1 0 25116 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_273
timestamp 1644511149
transform 1 0 26220 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_279
timestamp 1644511149
transform 1 0 26772 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_281
timestamp 1644511149
transform 1 0 26956 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_293
timestamp 1644511149
transform 1 0 28060 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_305
timestamp 1644511149
transform 1 0 29164 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_317
timestamp 1644511149
transform 1 0 30268 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_329
timestamp 1644511149
transform 1 0 31372 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_335
timestamp 1644511149
transform 1 0 31924 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_337
timestamp 1644511149
transform 1 0 32108 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_349
timestamp 1644511149
transform 1 0 33212 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_361
timestamp 1644511149
transform 1 0 34316 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_373
timestamp 1644511149
transform 1 0 35420 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_385
timestamp 1644511149
transform 1 0 36524 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_391
timestamp 1644511149
transform 1 0 37076 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_393
timestamp 1644511149
transform 1 0 37260 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_405
timestamp 1644511149
transform 1 0 38364 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_417
timestamp 1644511149
transform 1 0 39468 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_429
timestamp 1644511149
transform 1 0 40572 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_441
timestamp 1644511149
transform 1 0 41676 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_447
timestamp 1644511149
transform 1 0 42228 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_449
timestamp 1644511149
transform 1 0 42412 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_461
timestamp 1644511149
transform 1 0 43516 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_473
timestamp 1644511149
transform 1 0 44620 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_485
timestamp 1644511149
transform 1 0 45724 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_497
timestamp 1644511149
transform 1 0 46828 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_503
timestamp 1644511149
transform 1 0 47380 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_505
timestamp 1644511149
transform 1 0 47564 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_517
timestamp 1644511149
transform 1 0 48668 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_529
timestamp 1644511149
transform 1 0 49772 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_541
timestamp 1644511149
transform 1 0 50876 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_553
timestamp 1644511149
transform 1 0 51980 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_559
timestamp 1644511149
transform 1 0 52532 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_561
timestamp 1644511149
transform 1 0 52716 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_573
timestamp 1644511149
transform 1 0 53820 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_585
timestamp 1644511149
transform 1 0 54924 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_597
timestamp 1644511149
transform 1 0 56028 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_609
timestamp 1644511149
transform 1 0 57132 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_615
timestamp 1644511149
transform 1 0 57684 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_617
timestamp 1644511149
transform 1 0 57868 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_629
timestamp 1644511149
transform 1 0 58972 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_641
timestamp 1644511149
transform 1 0 60076 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_653
timestamp 1644511149
transform 1 0 61180 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_665
timestamp 1644511149
transform 1 0 62284 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_671
timestamp 1644511149
transform 1 0 62836 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_673
timestamp 1644511149
transform 1 0 63020 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_685
timestamp 1644511149
transform 1 0 64124 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_697
timestamp 1644511149
transform 1 0 65228 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_709
timestamp 1644511149
transform 1 0 66332 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_721
timestamp 1644511149
transform 1 0 67436 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_727
timestamp 1644511149
transform 1 0 67988 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_729
timestamp 1644511149
transform 1 0 68172 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_741
timestamp 1644511149
transform 1 0 69276 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_753
timestamp 1644511149
transform 1 0 70380 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_765
timestamp 1644511149
transform 1 0 71484 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_777
timestamp 1644511149
transform 1 0 72588 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_783
timestamp 1644511149
transform 1 0 73140 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_785
timestamp 1644511149
transform 1 0 73324 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_797
timestamp 1644511149
transform 1 0 74428 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_809
timestamp 1644511149
transform 1 0 75532 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_821
timestamp 1644511149
transform 1 0 76636 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_827
timestamp 1644511149
transform 1 0 77188 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_41_830
timestamp 1644511149
transform 1 0 77464 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_836
timestamp 1644511149
transform 1 0 78016 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_841
timestamp 1644511149
transform 1 0 78476 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_3
timestamp 1644511149
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_15
timestamp 1644511149
transform 1 0 2484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_27
timestamp 1644511149
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_29
timestamp 1644511149
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_41
timestamp 1644511149
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_53
timestamp 1644511149
transform 1 0 5980 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_65
timestamp 1644511149
transform 1 0 7084 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_77
timestamp 1644511149
transform 1 0 8188 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_83
timestamp 1644511149
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_85
timestamp 1644511149
transform 1 0 8924 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_97
timestamp 1644511149
transform 1 0 10028 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_109
timestamp 1644511149
transform 1 0 11132 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_121
timestamp 1644511149
transform 1 0 12236 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_133
timestamp 1644511149
transform 1 0 13340 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_139
timestamp 1644511149
transform 1 0 13892 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_141
timestamp 1644511149
transform 1 0 14076 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_153
timestamp 1644511149
transform 1 0 15180 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_165
timestamp 1644511149
transform 1 0 16284 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_177
timestamp 1644511149
transform 1 0 17388 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_189
timestamp 1644511149
transform 1 0 18492 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_195
timestamp 1644511149
transform 1 0 19044 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_197
timestamp 1644511149
transform 1 0 19228 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_209
timestamp 1644511149
transform 1 0 20332 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_221
timestamp 1644511149
transform 1 0 21436 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_233
timestamp 1644511149
transform 1 0 22540 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_245
timestamp 1644511149
transform 1 0 23644 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_251
timestamp 1644511149
transform 1 0 24196 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_253
timestamp 1644511149
transform 1 0 24380 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_265
timestamp 1644511149
transform 1 0 25484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_277
timestamp 1644511149
transform 1 0 26588 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_289
timestamp 1644511149
transform 1 0 27692 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_301
timestamp 1644511149
transform 1 0 28796 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_307
timestamp 1644511149
transform 1 0 29348 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_309
timestamp 1644511149
transform 1 0 29532 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_321
timestamp 1644511149
transform 1 0 30636 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_333
timestamp 1644511149
transform 1 0 31740 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_345
timestamp 1644511149
transform 1 0 32844 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_357
timestamp 1644511149
transform 1 0 33948 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_363
timestamp 1644511149
transform 1 0 34500 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_365
timestamp 1644511149
transform 1 0 34684 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_377
timestamp 1644511149
transform 1 0 35788 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_389
timestamp 1644511149
transform 1 0 36892 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_401
timestamp 1644511149
transform 1 0 37996 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_413
timestamp 1644511149
transform 1 0 39100 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_419
timestamp 1644511149
transform 1 0 39652 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_421
timestamp 1644511149
transform 1 0 39836 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_433
timestamp 1644511149
transform 1 0 40940 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_445
timestamp 1644511149
transform 1 0 42044 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_457
timestamp 1644511149
transform 1 0 43148 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_469
timestamp 1644511149
transform 1 0 44252 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_475
timestamp 1644511149
transform 1 0 44804 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_477
timestamp 1644511149
transform 1 0 44988 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_489
timestamp 1644511149
transform 1 0 46092 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_501
timestamp 1644511149
transform 1 0 47196 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_513
timestamp 1644511149
transform 1 0 48300 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_525
timestamp 1644511149
transform 1 0 49404 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_531
timestamp 1644511149
transform 1 0 49956 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_533
timestamp 1644511149
transform 1 0 50140 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_545
timestamp 1644511149
transform 1 0 51244 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_557
timestamp 1644511149
transform 1 0 52348 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_569
timestamp 1644511149
transform 1 0 53452 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_581
timestamp 1644511149
transform 1 0 54556 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_587
timestamp 1644511149
transform 1 0 55108 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_589
timestamp 1644511149
transform 1 0 55292 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_601
timestamp 1644511149
transform 1 0 56396 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_613
timestamp 1644511149
transform 1 0 57500 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_625
timestamp 1644511149
transform 1 0 58604 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_637
timestamp 1644511149
transform 1 0 59708 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_643
timestamp 1644511149
transform 1 0 60260 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_645
timestamp 1644511149
transform 1 0 60444 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_657
timestamp 1644511149
transform 1 0 61548 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_669
timestamp 1644511149
transform 1 0 62652 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_681
timestamp 1644511149
transform 1 0 63756 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_693
timestamp 1644511149
transform 1 0 64860 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_699
timestamp 1644511149
transform 1 0 65412 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_701
timestamp 1644511149
transform 1 0 65596 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_713
timestamp 1644511149
transform 1 0 66700 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_725
timestamp 1644511149
transform 1 0 67804 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_737
timestamp 1644511149
transform 1 0 68908 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_749
timestamp 1644511149
transform 1 0 70012 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_755
timestamp 1644511149
transform 1 0 70564 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_757
timestamp 1644511149
transform 1 0 70748 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_769
timestamp 1644511149
transform 1 0 71852 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_781
timestamp 1644511149
transform 1 0 72956 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_793
timestamp 1644511149
transform 1 0 74060 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_805
timestamp 1644511149
transform 1 0 75164 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_811
timestamp 1644511149
transform 1 0 75716 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_813
timestamp 1644511149
transform 1 0 75900 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_825
timestamp 1644511149
transform 1 0 77004 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_837
timestamp 1644511149
transform 1 0 78108 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_841
timestamp 1644511149
transform 1 0 78476 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_3
timestamp 1644511149
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_15
timestamp 1644511149
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_27
timestamp 1644511149
transform 1 0 3588 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_39
timestamp 1644511149
transform 1 0 4692 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_51
timestamp 1644511149
transform 1 0 5796 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_55
timestamp 1644511149
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_57
timestamp 1644511149
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_69
timestamp 1644511149
transform 1 0 7452 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_81
timestamp 1644511149
transform 1 0 8556 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_93
timestamp 1644511149
transform 1 0 9660 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_105
timestamp 1644511149
transform 1 0 10764 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_111
timestamp 1644511149
transform 1 0 11316 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_113
timestamp 1644511149
transform 1 0 11500 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_125
timestamp 1644511149
transform 1 0 12604 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_137
timestamp 1644511149
transform 1 0 13708 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_149
timestamp 1644511149
transform 1 0 14812 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_161
timestamp 1644511149
transform 1 0 15916 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_167
timestamp 1644511149
transform 1 0 16468 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_169
timestamp 1644511149
transform 1 0 16652 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_181
timestamp 1644511149
transform 1 0 17756 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_193
timestamp 1644511149
transform 1 0 18860 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_205
timestamp 1644511149
transform 1 0 19964 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_217
timestamp 1644511149
transform 1 0 21068 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_223
timestamp 1644511149
transform 1 0 21620 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_225
timestamp 1644511149
transform 1 0 21804 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_237
timestamp 1644511149
transform 1 0 22908 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_249
timestamp 1644511149
transform 1 0 24012 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_261
timestamp 1644511149
transform 1 0 25116 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_273
timestamp 1644511149
transform 1 0 26220 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_279
timestamp 1644511149
transform 1 0 26772 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_281
timestamp 1644511149
transform 1 0 26956 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_293
timestamp 1644511149
transform 1 0 28060 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_305
timestamp 1644511149
transform 1 0 29164 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_317
timestamp 1644511149
transform 1 0 30268 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_329
timestamp 1644511149
transform 1 0 31372 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_335
timestamp 1644511149
transform 1 0 31924 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_337
timestamp 1644511149
transform 1 0 32108 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_349
timestamp 1644511149
transform 1 0 33212 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_361
timestamp 1644511149
transform 1 0 34316 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_373
timestamp 1644511149
transform 1 0 35420 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_385
timestamp 1644511149
transform 1 0 36524 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_391
timestamp 1644511149
transform 1 0 37076 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_393
timestamp 1644511149
transform 1 0 37260 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_405
timestamp 1644511149
transform 1 0 38364 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_43_419
timestamp 1644511149
transform 1 0 39652 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_43_427
timestamp 1644511149
transform 1 0 40388 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_439
timestamp 1644511149
transform 1 0 41492 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_447
timestamp 1644511149
transform 1 0 42228 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_449
timestamp 1644511149
transform 1 0 42412 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_461
timestamp 1644511149
transform 1 0 43516 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_473
timestamp 1644511149
transform 1 0 44620 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_485
timestamp 1644511149
transform 1 0 45724 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_497
timestamp 1644511149
transform 1 0 46828 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_503
timestamp 1644511149
transform 1 0 47380 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_505
timestamp 1644511149
transform 1 0 47564 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_517
timestamp 1644511149
transform 1 0 48668 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_529
timestamp 1644511149
transform 1 0 49772 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_541
timestamp 1644511149
transform 1 0 50876 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_553
timestamp 1644511149
transform 1 0 51980 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_559
timestamp 1644511149
transform 1 0 52532 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_561
timestamp 1644511149
transform 1 0 52716 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_573
timestamp 1644511149
transform 1 0 53820 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_585
timestamp 1644511149
transform 1 0 54924 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_597
timestamp 1644511149
transform 1 0 56028 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_609
timestamp 1644511149
transform 1 0 57132 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_615
timestamp 1644511149
transform 1 0 57684 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_617
timestamp 1644511149
transform 1 0 57868 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_629
timestamp 1644511149
transform 1 0 58972 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_641
timestamp 1644511149
transform 1 0 60076 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_653
timestamp 1644511149
transform 1 0 61180 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_665
timestamp 1644511149
transform 1 0 62284 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_671
timestamp 1644511149
transform 1 0 62836 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_673
timestamp 1644511149
transform 1 0 63020 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_685
timestamp 1644511149
transform 1 0 64124 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_697
timestamp 1644511149
transform 1 0 65228 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_709
timestamp 1644511149
transform 1 0 66332 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_721
timestamp 1644511149
transform 1 0 67436 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_727
timestamp 1644511149
transform 1 0 67988 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_729
timestamp 1644511149
transform 1 0 68172 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_741
timestamp 1644511149
transform 1 0 69276 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_753
timestamp 1644511149
transform 1 0 70380 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_765
timestamp 1644511149
transform 1 0 71484 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_777
timestamp 1644511149
transform 1 0 72588 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_783
timestamp 1644511149
transform 1 0 73140 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_785
timestamp 1644511149
transform 1 0 73324 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_797
timestamp 1644511149
transform 1 0 74428 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_809
timestamp 1644511149
transform 1 0 75532 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_821
timestamp 1644511149
transform 1 0 76636 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_833
timestamp 1644511149
transform 1 0 77740 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_839
timestamp 1644511149
transform 1 0 78292 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_43_841
timestamp 1644511149
transform 1 0 78476 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_3
timestamp 1644511149
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_15
timestamp 1644511149
transform 1 0 2484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp 1644511149
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_29
timestamp 1644511149
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_41
timestamp 1644511149
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_53
timestamp 1644511149
transform 1 0 5980 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_65
timestamp 1644511149
transform 1 0 7084 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_77
timestamp 1644511149
transform 1 0 8188 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_83
timestamp 1644511149
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_85
timestamp 1644511149
transform 1 0 8924 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_97
timestamp 1644511149
transform 1 0 10028 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_109
timestamp 1644511149
transform 1 0 11132 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_121
timestamp 1644511149
transform 1 0 12236 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_133
timestamp 1644511149
transform 1 0 13340 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_139
timestamp 1644511149
transform 1 0 13892 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_141
timestamp 1644511149
transform 1 0 14076 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_153
timestamp 1644511149
transform 1 0 15180 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_165
timestamp 1644511149
transform 1 0 16284 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_177
timestamp 1644511149
transform 1 0 17388 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_189
timestamp 1644511149
transform 1 0 18492 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_195
timestamp 1644511149
transform 1 0 19044 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_197
timestamp 1644511149
transform 1 0 19228 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_209
timestamp 1644511149
transform 1 0 20332 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_221
timestamp 1644511149
transform 1 0 21436 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_233
timestamp 1644511149
transform 1 0 22540 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_245
timestamp 1644511149
transform 1 0 23644 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_251
timestamp 1644511149
transform 1 0 24196 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_253
timestamp 1644511149
transform 1 0 24380 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_265
timestamp 1644511149
transform 1 0 25484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_277
timestamp 1644511149
transform 1 0 26588 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_289
timestamp 1644511149
transform 1 0 27692 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_301
timestamp 1644511149
transform 1 0 28796 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_307
timestamp 1644511149
transform 1 0 29348 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_309
timestamp 1644511149
transform 1 0 29532 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_321
timestamp 1644511149
transform 1 0 30636 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_333
timestamp 1644511149
transform 1 0 31740 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_345
timestamp 1644511149
transform 1 0 32844 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_357
timestamp 1644511149
transform 1 0 33948 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_363
timestamp 1644511149
transform 1 0 34500 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_365
timestamp 1644511149
transform 1 0 34684 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_377
timestamp 1644511149
transform 1 0 35788 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_389
timestamp 1644511149
transform 1 0 36892 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_401
timestamp 1644511149
transform 1 0 37996 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_413
timestamp 1644511149
transform 1 0 39100 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_419
timestamp 1644511149
transform 1 0 39652 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_421
timestamp 1644511149
transform 1 0 39836 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_433
timestamp 1644511149
transform 1 0 40940 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_445
timestamp 1644511149
transform 1 0 42044 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_457
timestamp 1644511149
transform 1 0 43148 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_469
timestamp 1644511149
transform 1 0 44252 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_475
timestamp 1644511149
transform 1 0 44804 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_477
timestamp 1644511149
transform 1 0 44988 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_489
timestamp 1644511149
transform 1 0 46092 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_501
timestamp 1644511149
transform 1 0 47196 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_513
timestamp 1644511149
transform 1 0 48300 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_525
timestamp 1644511149
transform 1 0 49404 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_531
timestamp 1644511149
transform 1 0 49956 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_533
timestamp 1644511149
transform 1 0 50140 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_545
timestamp 1644511149
transform 1 0 51244 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_557
timestamp 1644511149
transform 1 0 52348 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_569
timestamp 1644511149
transform 1 0 53452 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_581
timestamp 1644511149
transform 1 0 54556 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_587
timestamp 1644511149
transform 1 0 55108 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_589
timestamp 1644511149
transform 1 0 55292 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_601
timestamp 1644511149
transform 1 0 56396 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_613
timestamp 1644511149
transform 1 0 57500 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_625
timestamp 1644511149
transform 1 0 58604 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_637
timestamp 1644511149
transform 1 0 59708 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_643
timestamp 1644511149
transform 1 0 60260 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_645
timestamp 1644511149
transform 1 0 60444 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_657
timestamp 1644511149
transform 1 0 61548 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_669
timestamp 1644511149
transform 1 0 62652 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_681
timestamp 1644511149
transform 1 0 63756 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_693
timestamp 1644511149
transform 1 0 64860 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_699
timestamp 1644511149
transform 1 0 65412 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_701
timestamp 1644511149
transform 1 0 65596 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_713
timestamp 1644511149
transform 1 0 66700 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_725
timestamp 1644511149
transform 1 0 67804 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_737
timestamp 1644511149
transform 1 0 68908 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_749
timestamp 1644511149
transform 1 0 70012 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_755
timestamp 1644511149
transform 1 0 70564 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_757
timestamp 1644511149
transform 1 0 70748 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_769
timestamp 1644511149
transform 1 0 71852 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_781
timestamp 1644511149
transform 1 0 72956 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_793
timestamp 1644511149
transform 1 0 74060 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_805
timestamp 1644511149
transform 1 0 75164 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_811
timestamp 1644511149
transform 1 0 75716 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_813
timestamp 1644511149
transform 1 0 75900 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_825
timestamp 1644511149
transform 1 0 77004 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_837
timestamp 1644511149
transform 1 0 78108 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_841
timestamp 1644511149
transform 1 0 78476 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_3
timestamp 1644511149
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_15
timestamp 1644511149
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_27
timestamp 1644511149
transform 1 0 3588 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_39
timestamp 1644511149
transform 1 0 4692 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_51
timestamp 1644511149
transform 1 0 5796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_55
timestamp 1644511149
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_57
timestamp 1644511149
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_69
timestamp 1644511149
transform 1 0 7452 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_81
timestamp 1644511149
transform 1 0 8556 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_93
timestamp 1644511149
transform 1 0 9660 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_105
timestamp 1644511149
transform 1 0 10764 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_111
timestamp 1644511149
transform 1 0 11316 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_113
timestamp 1644511149
transform 1 0 11500 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_125
timestamp 1644511149
transform 1 0 12604 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_137
timestamp 1644511149
transform 1 0 13708 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_149
timestamp 1644511149
transform 1 0 14812 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_161
timestamp 1644511149
transform 1 0 15916 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_167
timestamp 1644511149
transform 1 0 16468 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_169
timestamp 1644511149
transform 1 0 16652 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_181
timestamp 1644511149
transform 1 0 17756 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_193
timestamp 1644511149
transform 1 0 18860 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_205
timestamp 1644511149
transform 1 0 19964 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_217
timestamp 1644511149
transform 1 0 21068 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_223
timestamp 1644511149
transform 1 0 21620 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_225
timestamp 1644511149
transform 1 0 21804 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_237
timestamp 1644511149
transform 1 0 22908 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_249
timestamp 1644511149
transform 1 0 24012 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_261
timestamp 1644511149
transform 1 0 25116 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_273
timestamp 1644511149
transform 1 0 26220 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_279
timestamp 1644511149
transform 1 0 26772 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_281
timestamp 1644511149
transform 1 0 26956 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_293
timestamp 1644511149
transform 1 0 28060 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_305
timestamp 1644511149
transform 1 0 29164 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_317
timestamp 1644511149
transform 1 0 30268 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_329
timestamp 1644511149
transform 1 0 31372 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_335
timestamp 1644511149
transform 1 0 31924 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_337
timestamp 1644511149
transform 1 0 32108 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_349
timestamp 1644511149
transform 1 0 33212 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_361
timestamp 1644511149
transform 1 0 34316 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_373
timestamp 1644511149
transform 1 0 35420 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_385
timestamp 1644511149
transform 1 0 36524 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_391
timestamp 1644511149
transform 1 0 37076 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_393
timestamp 1644511149
transform 1 0 37260 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_405
timestamp 1644511149
transform 1 0 38364 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_417
timestamp 1644511149
transform 1 0 39468 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_429
timestamp 1644511149
transform 1 0 40572 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_441
timestamp 1644511149
transform 1 0 41676 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_447
timestamp 1644511149
transform 1 0 42228 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_449
timestamp 1644511149
transform 1 0 42412 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_461
timestamp 1644511149
transform 1 0 43516 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_473
timestamp 1644511149
transform 1 0 44620 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_485
timestamp 1644511149
transform 1 0 45724 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_497
timestamp 1644511149
transform 1 0 46828 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_503
timestamp 1644511149
transform 1 0 47380 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_505
timestamp 1644511149
transform 1 0 47564 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_517
timestamp 1644511149
transform 1 0 48668 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_529
timestamp 1644511149
transform 1 0 49772 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_541
timestamp 1644511149
transform 1 0 50876 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_553
timestamp 1644511149
transform 1 0 51980 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_559
timestamp 1644511149
transform 1 0 52532 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_561
timestamp 1644511149
transform 1 0 52716 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_573
timestamp 1644511149
transform 1 0 53820 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_585
timestamp 1644511149
transform 1 0 54924 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_597
timestamp 1644511149
transform 1 0 56028 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_609
timestamp 1644511149
transform 1 0 57132 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_615
timestamp 1644511149
transform 1 0 57684 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_617
timestamp 1644511149
transform 1 0 57868 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_629
timestamp 1644511149
transform 1 0 58972 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_641
timestamp 1644511149
transform 1 0 60076 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_653
timestamp 1644511149
transform 1 0 61180 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_665
timestamp 1644511149
transform 1 0 62284 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_671
timestamp 1644511149
transform 1 0 62836 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_673
timestamp 1644511149
transform 1 0 63020 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_685
timestamp 1644511149
transform 1 0 64124 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_697
timestamp 1644511149
transform 1 0 65228 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_709
timestamp 1644511149
transform 1 0 66332 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_721
timestamp 1644511149
transform 1 0 67436 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_727
timestamp 1644511149
transform 1 0 67988 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_729
timestamp 1644511149
transform 1 0 68172 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_741
timestamp 1644511149
transform 1 0 69276 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_753
timestamp 1644511149
transform 1 0 70380 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_765
timestamp 1644511149
transform 1 0 71484 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_777
timestamp 1644511149
transform 1 0 72588 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_783
timestamp 1644511149
transform 1 0 73140 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_785
timestamp 1644511149
transform 1 0 73324 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_797
timestamp 1644511149
transform 1 0 74428 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_809
timestamp 1644511149
transform 1 0 75532 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_821
timestamp 1644511149
transform 1 0 76636 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_833
timestamp 1644511149
transform 1 0 77740 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_839
timestamp 1644511149
transform 1 0 78292 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_45_841
timestamp 1644511149
transform 1 0 78476 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_9
timestamp 1644511149
transform 1 0 1932 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_21
timestamp 1644511149
transform 1 0 3036 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_27
timestamp 1644511149
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_29
timestamp 1644511149
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_41
timestamp 1644511149
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_53
timestamp 1644511149
transform 1 0 5980 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_65
timestamp 1644511149
transform 1 0 7084 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_77
timestamp 1644511149
transform 1 0 8188 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_83
timestamp 1644511149
transform 1 0 8740 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_85
timestamp 1644511149
transform 1 0 8924 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_97
timestamp 1644511149
transform 1 0 10028 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_109
timestamp 1644511149
transform 1 0 11132 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_121
timestamp 1644511149
transform 1 0 12236 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_133
timestamp 1644511149
transform 1 0 13340 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_139
timestamp 1644511149
transform 1 0 13892 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_141
timestamp 1644511149
transform 1 0 14076 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_153
timestamp 1644511149
transform 1 0 15180 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_165
timestamp 1644511149
transform 1 0 16284 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_177
timestamp 1644511149
transform 1 0 17388 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_189
timestamp 1644511149
transform 1 0 18492 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_195
timestamp 1644511149
transform 1 0 19044 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_197
timestamp 1644511149
transform 1 0 19228 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_209
timestamp 1644511149
transform 1 0 20332 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_221
timestamp 1644511149
transform 1 0 21436 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_233
timestamp 1644511149
transform 1 0 22540 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_245
timestamp 1644511149
transform 1 0 23644 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_251
timestamp 1644511149
transform 1 0 24196 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_253
timestamp 1644511149
transform 1 0 24380 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_265
timestamp 1644511149
transform 1 0 25484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_277
timestamp 1644511149
transform 1 0 26588 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_289
timestamp 1644511149
transform 1 0 27692 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_301
timestamp 1644511149
transform 1 0 28796 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_307
timestamp 1644511149
transform 1 0 29348 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_309
timestamp 1644511149
transform 1 0 29532 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_321
timestamp 1644511149
transform 1 0 30636 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_333
timestamp 1644511149
transform 1 0 31740 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_345
timestamp 1644511149
transform 1 0 32844 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_357
timestamp 1644511149
transform 1 0 33948 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_363
timestamp 1644511149
transform 1 0 34500 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_365
timestamp 1644511149
transform 1 0 34684 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_377
timestamp 1644511149
transform 1 0 35788 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_389
timestamp 1644511149
transform 1 0 36892 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_401
timestamp 1644511149
transform 1 0 37996 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_413
timestamp 1644511149
transform 1 0 39100 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_419
timestamp 1644511149
transform 1 0 39652 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_421
timestamp 1644511149
transform 1 0 39836 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_433
timestamp 1644511149
transform 1 0 40940 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_445
timestamp 1644511149
transform 1 0 42044 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_457
timestamp 1644511149
transform 1 0 43148 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_469
timestamp 1644511149
transform 1 0 44252 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_475
timestamp 1644511149
transform 1 0 44804 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_477
timestamp 1644511149
transform 1 0 44988 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_489
timestamp 1644511149
transform 1 0 46092 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_501
timestamp 1644511149
transform 1 0 47196 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_513
timestamp 1644511149
transform 1 0 48300 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_525
timestamp 1644511149
transform 1 0 49404 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_531
timestamp 1644511149
transform 1 0 49956 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_533
timestamp 1644511149
transform 1 0 50140 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_545
timestamp 1644511149
transform 1 0 51244 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_557
timestamp 1644511149
transform 1 0 52348 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_569
timestamp 1644511149
transform 1 0 53452 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_581
timestamp 1644511149
transform 1 0 54556 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_587
timestamp 1644511149
transform 1 0 55108 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_589
timestamp 1644511149
transform 1 0 55292 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_601
timestamp 1644511149
transform 1 0 56396 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_613
timestamp 1644511149
transform 1 0 57500 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_625
timestamp 1644511149
transform 1 0 58604 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_637
timestamp 1644511149
transform 1 0 59708 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_643
timestamp 1644511149
transform 1 0 60260 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_645
timestamp 1644511149
transform 1 0 60444 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_657
timestamp 1644511149
transform 1 0 61548 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_669
timestamp 1644511149
transform 1 0 62652 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_681
timestamp 1644511149
transform 1 0 63756 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_693
timestamp 1644511149
transform 1 0 64860 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_699
timestamp 1644511149
transform 1 0 65412 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_701
timestamp 1644511149
transform 1 0 65596 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_713
timestamp 1644511149
transform 1 0 66700 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_725
timestamp 1644511149
transform 1 0 67804 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_737
timestamp 1644511149
transform 1 0 68908 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_749
timestamp 1644511149
transform 1 0 70012 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_755
timestamp 1644511149
transform 1 0 70564 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_757
timestamp 1644511149
transform 1 0 70748 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_769
timestamp 1644511149
transform 1 0 71852 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_781
timestamp 1644511149
transform 1 0 72956 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_793
timestamp 1644511149
transform 1 0 74060 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_805
timestamp 1644511149
transform 1 0 75164 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_811
timestamp 1644511149
transform 1 0 75716 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_813
timestamp 1644511149
transform 1 0 75900 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_825
timestamp 1644511149
transform 1 0 77004 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_837
timestamp 1644511149
transform 1 0 78108 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_841
timestamp 1644511149
transform 1 0 78476 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_3
timestamp 1644511149
transform 1 0 1380 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_15
timestamp 1644511149
transform 1 0 2484 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_27
timestamp 1644511149
transform 1 0 3588 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_39
timestamp 1644511149
transform 1 0 4692 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_51
timestamp 1644511149
transform 1 0 5796 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_55
timestamp 1644511149
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_57
timestamp 1644511149
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_69
timestamp 1644511149
transform 1 0 7452 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_81
timestamp 1644511149
transform 1 0 8556 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_93
timestamp 1644511149
transform 1 0 9660 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_105
timestamp 1644511149
transform 1 0 10764 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_111
timestamp 1644511149
transform 1 0 11316 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_113
timestamp 1644511149
transform 1 0 11500 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_125
timestamp 1644511149
transform 1 0 12604 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_137
timestamp 1644511149
transform 1 0 13708 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_149
timestamp 1644511149
transform 1 0 14812 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_161
timestamp 1644511149
transform 1 0 15916 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_167
timestamp 1644511149
transform 1 0 16468 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_169
timestamp 1644511149
transform 1 0 16652 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_181
timestamp 1644511149
transform 1 0 17756 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_193
timestamp 1644511149
transform 1 0 18860 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_205
timestamp 1644511149
transform 1 0 19964 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_217
timestamp 1644511149
transform 1 0 21068 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_223
timestamp 1644511149
transform 1 0 21620 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_225
timestamp 1644511149
transform 1 0 21804 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_237
timestamp 1644511149
transform 1 0 22908 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_249
timestamp 1644511149
transform 1 0 24012 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_261
timestamp 1644511149
transform 1 0 25116 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_273
timestamp 1644511149
transform 1 0 26220 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_279
timestamp 1644511149
transform 1 0 26772 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_281
timestamp 1644511149
transform 1 0 26956 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_293
timestamp 1644511149
transform 1 0 28060 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_305
timestamp 1644511149
transform 1 0 29164 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_317
timestamp 1644511149
transform 1 0 30268 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_329
timestamp 1644511149
transform 1 0 31372 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_335
timestamp 1644511149
transform 1 0 31924 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_337
timestamp 1644511149
transform 1 0 32108 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_349
timestamp 1644511149
transform 1 0 33212 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_361
timestamp 1644511149
transform 1 0 34316 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_373
timestamp 1644511149
transform 1 0 35420 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_385
timestamp 1644511149
transform 1 0 36524 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_391
timestamp 1644511149
transform 1 0 37076 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_393
timestamp 1644511149
transform 1 0 37260 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_405
timestamp 1644511149
transform 1 0 38364 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_417
timestamp 1644511149
transform 1 0 39468 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_429
timestamp 1644511149
transform 1 0 40572 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_441
timestamp 1644511149
transform 1 0 41676 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_447
timestamp 1644511149
transform 1 0 42228 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_449
timestamp 1644511149
transform 1 0 42412 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_461
timestamp 1644511149
transform 1 0 43516 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_473
timestamp 1644511149
transform 1 0 44620 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_485
timestamp 1644511149
transform 1 0 45724 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_497
timestamp 1644511149
transform 1 0 46828 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_503
timestamp 1644511149
transform 1 0 47380 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_505
timestamp 1644511149
transform 1 0 47564 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_517
timestamp 1644511149
transform 1 0 48668 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_529
timestamp 1644511149
transform 1 0 49772 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_541
timestamp 1644511149
transform 1 0 50876 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_553
timestamp 1644511149
transform 1 0 51980 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_559
timestamp 1644511149
transform 1 0 52532 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_561
timestamp 1644511149
transform 1 0 52716 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_573
timestamp 1644511149
transform 1 0 53820 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_585
timestamp 1644511149
transform 1 0 54924 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_597
timestamp 1644511149
transform 1 0 56028 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_609
timestamp 1644511149
transform 1 0 57132 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_615
timestamp 1644511149
transform 1 0 57684 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_617
timestamp 1644511149
transform 1 0 57868 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_629
timestamp 1644511149
transform 1 0 58972 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_641
timestamp 1644511149
transform 1 0 60076 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_653
timestamp 1644511149
transform 1 0 61180 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_665
timestamp 1644511149
transform 1 0 62284 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_671
timestamp 1644511149
transform 1 0 62836 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_673
timestamp 1644511149
transform 1 0 63020 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_685
timestamp 1644511149
transform 1 0 64124 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_697
timestamp 1644511149
transform 1 0 65228 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_709
timestamp 1644511149
transform 1 0 66332 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_721
timestamp 1644511149
transform 1 0 67436 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_727
timestamp 1644511149
transform 1 0 67988 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_729
timestamp 1644511149
transform 1 0 68172 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_741
timestamp 1644511149
transform 1 0 69276 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_753
timestamp 1644511149
transform 1 0 70380 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_765
timestamp 1644511149
transform 1 0 71484 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_777
timestamp 1644511149
transform 1 0 72588 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_783
timestamp 1644511149
transform 1 0 73140 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_785
timestamp 1644511149
transform 1 0 73324 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_797
timestamp 1644511149
transform 1 0 74428 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_809
timestamp 1644511149
transform 1 0 75532 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_821
timestamp 1644511149
transform 1 0 76636 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_836
timestamp 1644511149
transform 1 0 78016 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_841
timestamp 1644511149
transform 1 0 78476 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_3
timestamp 1644511149
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_15
timestamp 1644511149
transform 1 0 2484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 1644511149
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_29
timestamp 1644511149
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_41
timestamp 1644511149
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_53
timestamp 1644511149
transform 1 0 5980 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_65
timestamp 1644511149
transform 1 0 7084 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_77
timestamp 1644511149
transform 1 0 8188 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_83
timestamp 1644511149
transform 1 0 8740 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_85
timestamp 1644511149
transform 1 0 8924 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_97
timestamp 1644511149
transform 1 0 10028 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_109
timestamp 1644511149
transform 1 0 11132 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_121
timestamp 1644511149
transform 1 0 12236 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_133
timestamp 1644511149
transform 1 0 13340 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_139
timestamp 1644511149
transform 1 0 13892 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_141
timestamp 1644511149
transform 1 0 14076 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_153
timestamp 1644511149
transform 1 0 15180 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_165
timestamp 1644511149
transform 1 0 16284 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_177
timestamp 1644511149
transform 1 0 17388 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_189
timestamp 1644511149
transform 1 0 18492 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_195
timestamp 1644511149
transform 1 0 19044 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_197
timestamp 1644511149
transform 1 0 19228 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_209
timestamp 1644511149
transform 1 0 20332 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_221
timestamp 1644511149
transform 1 0 21436 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_233
timestamp 1644511149
transform 1 0 22540 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_245
timestamp 1644511149
transform 1 0 23644 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_251
timestamp 1644511149
transform 1 0 24196 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_253
timestamp 1644511149
transform 1 0 24380 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_265
timestamp 1644511149
transform 1 0 25484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_277
timestamp 1644511149
transform 1 0 26588 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_289
timestamp 1644511149
transform 1 0 27692 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_301
timestamp 1644511149
transform 1 0 28796 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_307
timestamp 1644511149
transform 1 0 29348 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_309
timestamp 1644511149
transform 1 0 29532 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_321
timestamp 1644511149
transform 1 0 30636 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_333
timestamp 1644511149
transform 1 0 31740 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_345
timestamp 1644511149
transform 1 0 32844 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_357
timestamp 1644511149
transform 1 0 33948 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_363
timestamp 1644511149
transform 1 0 34500 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_365
timestamp 1644511149
transform 1 0 34684 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_377
timestamp 1644511149
transform 1 0 35788 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_389
timestamp 1644511149
transform 1 0 36892 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_401
timestamp 1644511149
transform 1 0 37996 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_413
timestamp 1644511149
transform 1 0 39100 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_419
timestamp 1644511149
transform 1 0 39652 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_421
timestamp 1644511149
transform 1 0 39836 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_433
timestamp 1644511149
transform 1 0 40940 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_445
timestamp 1644511149
transform 1 0 42044 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_457
timestamp 1644511149
transform 1 0 43148 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_469
timestamp 1644511149
transform 1 0 44252 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_475
timestamp 1644511149
transform 1 0 44804 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_477
timestamp 1644511149
transform 1 0 44988 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_489
timestamp 1644511149
transform 1 0 46092 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_501
timestamp 1644511149
transform 1 0 47196 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_513
timestamp 1644511149
transform 1 0 48300 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_525
timestamp 1644511149
transform 1 0 49404 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_531
timestamp 1644511149
transform 1 0 49956 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_533
timestamp 1644511149
transform 1 0 50140 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_545
timestamp 1644511149
transform 1 0 51244 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_557
timestamp 1644511149
transform 1 0 52348 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_569
timestamp 1644511149
transform 1 0 53452 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_581
timestamp 1644511149
transform 1 0 54556 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_587
timestamp 1644511149
transform 1 0 55108 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_589
timestamp 1644511149
transform 1 0 55292 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_601
timestamp 1644511149
transform 1 0 56396 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_613
timestamp 1644511149
transform 1 0 57500 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_625
timestamp 1644511149
transform 1 0 58604 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_637
timestamp 1644511149
transform 1 0 59708 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_643
timestamp 1644511149
transform 1 0 60260 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_645
timestamp 1644511149
transform 1 0 60444 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_657
timestamp 1644511149
transform 1 0 61548 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_669
timestamp 1644511149
transform 1 0 62652 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_681
timestamp 1644511149
transform 1 0 63756 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_693
timestamp 1644511149
transform 1 0 64860 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_699
timestamp 1644511149
transform 1 0 65412 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_701
timestamp 1644511149
transform 1 0 65596 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_713
timestamp 1644511149
transform 1 0 66700 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_725
timestamp 1644511149
transform 1 0 67804 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_737
timestamp 1644511149
transform 1 0 68908 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_749
timestamp 1644511149
transform 1 0 70012 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_755
timestamp 1644511149
transform 1 0 70564 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_757
timestamp 1644511149
transform 1 0 70748 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_769
timestamp 1644511149
transform 1 0 71852 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_781
timestamp 1644511149
transform 1 0 72956 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_793
timestamp 1644511149
transform 1 0 74060 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_805
timestamp 1644511149
transform 1 0 75164 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_811
timestamp 1644511149
transform 1 0 75716 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_813
timestamp 1644511149
transform 1 0 75900 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_825
timestamp 1644511149
transform 1 0 77004 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_837
timestamp 1644511149
transform 1 0 78108 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_841
timestamp 1644511149
transform 1 0 78476 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_3
timestamp 1644511149
transform 1 0 1380 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_15
timestamp 1644511149
transform 1 0 2484 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_27
timestamp 1644511149
transform 1 0 3588 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_39
timestamp 1644511149
transform 1 0 4692 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_51
timestamp 1644511149
transform 1 0 5796 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_55
timestamp 1644511149
transform 1 0 6164 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_57
timestamp 1644511149
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_69
timestamp 1644511149
transform 1 0 7452 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_81
timestamp 1644511149
transform 1 0 8556 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_93
timestamp 1644511149
transform 1 0 9660 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_105
timestamp 1644511149
transform 1 0 10764 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_111
timestamp 1644511149
transform 1 0 11316 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_113
timestamp 1644511149
transform 1 0 11500 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_125
timestamp 1644511149
transform 1 0 12604 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_137
timestamp 1644511149
transform 1 0 13708 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_149
timestamp 1644511149
transform 1 0 14812 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_161
timestamp 1644511149
transform 1 0 15916 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_167
timestamp 1644511149
transform 1 0 16468 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_169
timestamp 1644511149
transform 1 0 16652 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_181
timestamp 1644511149
transform 1 0 17756 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_193
timestamp 1644511149
transform 1 0 18860 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_205
timestamp 1644511149
transform 1 0 19964 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_217
timestamp 1644511149
transform 1 0 21068 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_223
timestamp 1644511149
transform 1 0 21620 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_225
timestamp 1644511149
transform 1 0 21804 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_237
timestamp 1644511149
transform 1 0 22908 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_249
timestamp 1644511149
transform 1 0 24012 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_261
timestamp 1644511149
transform 1 0 25116 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_273
timestamp 1644511149
transform 1 0 26220 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_279
timestamp 1644511149
transform 1 0 26772 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_281
timestamp 1644511149
transform 1 0 26956 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_293
timestamp 1644511149
transform 1 0 28060 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_305
timestamp 1644511149
transform 1 0 29164 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_317
timestamp 1644511149
transform 1 0 30268 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_329
timestamp 1644511149
transform 1 0 31372 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_335
timestamp 1644511149
transform 1 0 31924 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_337
timestamp 1644511149
transform 1 0 32108 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_349
timestamp 1644511149
transform 1 0 33212 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_361
timestamp 1644511149
transform 1 0 34316 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_373
timestamp 1644511149
transform 1 0 35420 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_385
timestamp 1644511149
transform 1 0 36524 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_391
timestamp 1644511149
transform 1 0 37076 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_393
timestamp 1644511149
transform 1 0 37260 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_405
timestamp 1644511149
transform 1 0 38364 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_417
timestamp 1644511149
transform 1 0 39468 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_429
timestamp 1644511149
transform 1 0 40572 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_441
timestamp 1644511149
transform 1 0 41676 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_447
timestamp 1644511149
transform 1 0 42228 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_449
timestamp 1644511149
transform 1 0 42412 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_461
timestamp 1644511149
transform 1 0 43516 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_473
timestamp 1644511149
transform 1 0 44620 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_485
timestamp 1644511149
transform 1 0 45724 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_497
timestamp 1644511149
transform 1 0 46828 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_503
timestamp 1644511149
transform 1 0 47380 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_505
timestamp 1644511149
transform 1 0 47564 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_517
timestamp 1644511149
transform 1 0 48668 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_529
timestamp 1644511149
transform 1 0 49772 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_541
timestamp 1644511149
transform 1 0 50876 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_553
timestamp 1644511149
transform 1 0 51980 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_559
timestamp 1644511149
transform 1 0 52532 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_561
timestamp 1644511149
transform 1 0 52716 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_573
timestamp 1644511149
transform 1 0 53820 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_585
timestamp 1644511149
transform 1 0 54924 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_597
timestamp 1644511149
transform 1 0 56028 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_609
timestamp 1644511149
transform 1 0 57132 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_615
timestamp 1644511149
transform 1 0 57684 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_617
timestamp 1644511149
transform 1 0 57868 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_629
timestamp 1644511149
transform 1 0 58972 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_641
timestamp 1644511149
transform 1 0 60076 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_653
timestamp 1644511149
transform 1 0 61180 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_665
timestamp 1644511149
transform 1 0 62284 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_671
timestamp 1644511149
transform 1 0 62836 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_673
timestamp 1644511149
transform 1 0 63020 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_685
timestamp 1644511149
transform 1 0 64124 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_697
timestamp 1644511149
transform 1 0 65228 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_709
timestamp 1644511149
transform 1 0 66332 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_721
timestamp 1644511149
transform 1 0 67436 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_727
timestamp 1644511149
transform 1 0 67988 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_729
timestamp 1644511149
transform 1 0 68172 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_741
timestamp 1644511149
transform 1 0 69276 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_753
timestamp 1644511149
transform 1 0 70380 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_765
timestamp 1644511149
transform 1 0 71484 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_777
timestamp 1644511149
transform 1 0 72588 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_783
timestamp 1644511149
transform 1 0 73140 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_785
timestamp 1644511149
transform 1 0 73324 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_797
timestamp 1644511149
transform 1 0 74428 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_809
timestamp 1644511149
transform 1 0 75532 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_821
timestamp 1644511149
transform 1 0 76636 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_833
timestamp 1644511149
transform 1 0 77740 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_839
timestamp 1644511149
transform 1 0 78292 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_49_841
timestamp 1644511149
transform 1 0 78476 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_3
timestamp 1644511149
transform 1 0 1380 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_15
timestamp 1644511149
transform 1 0 2484 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_27
timestamp 1644511149
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_29
timestamp 1644511149
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_41
timestamp 1644511149
transform 1 0 4876 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_53
timestamp 1644511149
transform 1 0 5980 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_65
timestamp 1644511149
transform 1 0 7084 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_77
timestamp 1644511149
transform 1 0 8188 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_83
timestamp 1644511149
transform 1 0 8740 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_85
timestamp 1644511149
transform 1 0 8924 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_97
timestamp 1644511149
transform 1 0 10028 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_109
timestamp 1644511149
transform 1 0 11132 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_121
timestamp 1644511149
transform 1 0 12236 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_133
timestamp 1644511149
transform 1 0 13340 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_139
timestamp 1644511149
transform 1 0 13892 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_141
timestamp 1644511149
transform 1 0 14076 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_153
timestamp 1644511149
transform 1 0 15180 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_165
timestamp 1644511149
transform 1 0 16284 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_177
timestamp 1644511149
transform 1 0 17388 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_189
timestamp 1644511149
transform 1 0 18492 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_195
timestamp 1644511149
transform 1 0 19044 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_197
timestamp 1644511149
transform 1 0 19228 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_209
timestamp 1644511149
transform 1 0 20332 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_221
timestamp 1644511149
transform 1 0 21436 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_233
timestamp 1644511149
transform 1 0 22540 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_245
timestamp 1644511149
transform 1 0 23644 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_251
timestamp 1644511149
transform 1 0 24196 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_253
timestamp 1644511149
transform 1 0 24380 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_265
timestamp 1644511149
transform 1 0 25484 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_277
timestamp 1644511149
transform 1 0 26588 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_289
timestamp 1644511149
transform 1 0 27692 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_301
timestamp 1644511149
transform 1 0 28796 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_307
timestamp 1644511149
transform 1 0 29348 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_309
timestamp 1644511149
transform 1 0 29532 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_321
timestamp 1644511149
transform 1 0 30636 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_333
timestamp 1644511149
transform 1 0 31740 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_345
timestamp 1644511149
transform 1 0 32844 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_357
timestamp 1644511149
transform 1 0 33948 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_363
timestamp 1644511149
transform 1 0 34500 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_365
timestamp 1644511149
transform 1 0 34684 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_377
timestamp 1644511149
transform 1 0 35788 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_389
timestamp 1644511149
transform 1 0 36892 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_401
timestamp 1644511149
transform 1 0 37996 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_413
timestamp 1644511149
transform 1 0 39100 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_419
timestamp 1644511149
transform 1 0 39652 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_421
timestamp 1644511149
transform 1 0 39836 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_433
timestamp 1644511149
transform 1 0 40940 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_445
timestamp 1644511149
transform 1 0 42044 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_457
timestamp 1644511149
transform 1 0 43148 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_469
timestamp 1644511149
transform 1 0 44252 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_475
timestamp 1644511149
transform 1 0 44804 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_477
timestamp 1644511149
transform 1 0 44988 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_489
timestamp 1644511149
transform 1 0 46092 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_501
timestamp 1644511149
transform 1 0 47196 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_513
timestamp 1644511149
transform 1 0 48300 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_525
timestamp 1644511149
transform 1 0 49404 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_531
timestamp 1644511149
transform 1 0 49956 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_533
timestamp 1644511149
transform 1 0 50140 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_545
timestamp 1644511149
transform 1 0 51244 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_557
timestamp 1644511149
transform 1 0 52348 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_569
timestamp 1644511149
transform 1 0 53452 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_581
timestamp 1644511149
transform 1 0 54556 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_587
timestamp 1644511149
transform 1 0 55108 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_589
timestamp 1644511149
transform 1 0 55292 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_601
timestamp 1644511149
transform 1 0 56396 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_613
timestamp 1644511149
transform 1 0 57500 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_625
timestamp 1644511149
transform 1 0 58604 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_637
timestamp 1644511149
transform 1 0 59708 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_643
timestamp 1644511149
transform 1 0 60260 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_645
timestamp 1644511149
transform 1 0 60444 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_657
timestamp 1644511149
transform 1 0 61548 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_669
timestamp 1644511149
transform 1 0 62652 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_681
timestamp 1644511149
transform 1 0 63756 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_693
timestamp 1644511149
transform 1 0 64860 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_699
timestamp 1644511149
transform 1 0 65412 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_701
timestamp 1644511149
transform 1 0 65596 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_713
timestamp 1644511149
transform 1 0 66700 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_725
timestamp 1644511149
transform 1 0 67804 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_737
timestamp 1644511149
transform 1 0 68908 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_749
timestamp 1644511149
transform 1 0 70012 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_755
timestamp 1644511149
transform 1 0 70564 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_757
timestamp 1644511149
transform 1 0 70748 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_769
timestamp 1644511149
transform 1 0 71852 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_781
timestamp 1644511149
transform 1 0 72956 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_793
timestamp 1644511149
transform 1 0 74060 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_805
timestamp 1644511149
transform 1 0 75164 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_811
timestamp 1644511149
transform 1 0 75716 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_813
timestamp 1644511149
transform 1 0 75900 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_825
timestamp 1644511149
transform 1 0 77004 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_837
timestamp 1644511149
transform 1 0 78108 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_841
timestamp 1644511149
transform 1 0 78476 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_3
timestamp 1644511149
transform 1 0 1380 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_15
timestamp 1644511149
transform 1 0 2484 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_27
timestamp 1644511149
transform 1 0 3588 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_39
timestamp 1644511149
transform 1 0 4692 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_51
timestamp 1644511149
transform 1 0 5796 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_55
timestamp 1644511149
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_57
timestamp 1644511149
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_69
timestamp 1644511149
transform 1 0 7452 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_81
timestamp 1644511149
transform 1 0 8556 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_93
timestamp 1644511149
transform 1 0 9660 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_105
timestamp 1644511149
transform 1 0 10764 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_111
timestamp 1644511149
transform 1 0 11316 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_113
timestamp 1644511149
transform 1 0 11500 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_125
timestamp 1644511149
transform 1 0 12604 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_137
timestamp 1644511149
transform 1 0 13708 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_149
timestamp 1644511149
transform 1 0 14812 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_161
timestamp 1644511149
transform 1 0 15916 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_167
timestamp 1644511149
transform 1 0 16468 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_169
timestamp 1644511149
transform 1 0 16652 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_181
timestamp 1644511149
transform 1 0 17756 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_193
timestamp 1644511149
transform 1 0 18860 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_205
timestamp 1644511149
transform 1 0 19964 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_217
timestamp 1644511149
transform 1 0 21068 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_223
timestamp 1644511149
transform 1 0 21620 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_225
timestamp 1644511149
transform 1 0 21804 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_237
timestamp 1644511149
transform 1 0 22908 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_249
timestamp 1644511149
transform 1 0 24012 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_261
timestamp 1644511149
transform 1 0 25116 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_273
timestamp 1644511149
transform 1 0 26220 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_279
timestamp 1644511149
transform 1 0 26772 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_281
timestamp 1644511149
transform 1 0 26956 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_293
timestamp 1644511149
transform 1 0 28060 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_305
timestamp 1644511149
transform 1 0 29164 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_317
timestamp 1644511149
transform 1 0 30268 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_329
timestamp 1644511149
transform 1 0 31372 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_335
timestamp 1644511149
transform 1 0 31924 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_337
timestamp 1644511149
transform 1 0 32108 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_349
timestamp 1644511149
transform 1 0 33212 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_361
timestamp 1644511149
transform 1 0 34316 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_373
timestamp 1644511149
transform 1 0 35420 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_385
timestamp 1644511149
transform 1 0 36524 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_391
timestamp 1644511149
transform 1 0 37076 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_393
timestamp 1644511149
transform 1 0 37260 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_405
timestamp 1644511149
transform 1 0 38364 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_417
timestamp 1644511149
transform 1 0 39468 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_429
timestamp 1644511149
transform 1 0 40572 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_441
timestamp 1644511149
transform 1 0 41676 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_447
timestamp 1644511149
transform 1 0 42228 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_449
timestamp 1644511149
transform 1 0 42412 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_461
timestamp 1644511149
transform 1 0 43516 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_473
timestamp 1644511149
transform 1 0 44620 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_485
timestamp 1644511149
transform 1 0 45724 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_497
timestamp 1644511149
transform 1 0 46828 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_503
timestamp 1644511149
transform 1 0 47380 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_505
timestamp 1644511149
transform 1 0 47564 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_517
timestamp 1644511149
transform 1 0 48668 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_529
timestamp 1644511149
transform 1 0 49772 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_541
timestamp 1644511149
transform 1 0 50876 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_553
timestamp 1644511149
transform 1 0 51980 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_559
timestamp 1644511149
transform 1 0 52532 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_561
timestamp 1644511149
transform 1 0 52716 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_573
timestamp 1644511149
transform 1 0 53820 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_585
timestamp 1644511149
transform 1 0 54924 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_597
timestamp 1644511149
transform 1 0 56028 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_609
timestamp 1644511149
transform 1 0 57132 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_615
timestamp 1644511149
transform 1 0 57684 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_617
timestamp 1644511149
transform 1 0 57868 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_629
timestamp 1644511149
transform 1 0 58972 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_641
timestamp 1644511149
transform 1 0 60076 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_653
timestamp 1644511149
transform 1 0 61180 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_665
timestamp 1644511149
transform 1 0 62284 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_671
timestamp 1644511149
transform 1 0 62836 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_673
timestamp 1644511149
transform 1 0 63020 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_685
timestamp 1644511149
transform 1 0 64124 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_697
timestamp 1644511149
transform 1 0 65228 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_709
timestamp 1644511149
transform 1 0 66332 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_721
timestamp 1644511149
transform 1 0 67436 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_727
timestamp 1644511149
transform 1 0 67988 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_729
timestamp 1644511149
transform 1 0 68172 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_741
timestamp 1644511149
transform 1 0 69276 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_753
timestamp 1644511149
transform 1 0 70380 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_765
timestamp 1644511149
transform 1 0 71484 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_777
timestamp 1644511149
transform 1 0 72588 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_783
timestamp 1644511149
transform 1 0 73140 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_785
timestamp 1644511149
transform 1 0 73324 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_797
timestamp 1644511149
transform 1 0 74428 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_809
timestamp 1644511149
transform 1 0 75532 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_821
timestamp 1644511149
transform 1 0 76636 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_833
timestamp 1644511149
transform 1 0 77740 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_839
timestamp 1644511149
transform 1 0 78292 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_51_841
timestamp 1644511149
transform 1 0 78476 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_3
timestamp 1644511149
transform 1 0 1380 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_15
timestamp 1644511149
transform 1 0 2484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_27
timestamp 1644511149
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_29
timestamp 1644511149
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_41
timestamp 1644511149
transform 1 0 4876 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_53
timestamp 1644511149
transform 1 0 5980 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_65
timestamp 1644511149
transform 1 0 7084 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_77
timestamp 1644511149
transform 1 0 8188 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_83
timestamp 1644511149
transform 1 0 8740 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_85
timestamp 1644511149
transform 1 0 8924 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_97
timestamp 1644511149
transform 1 0 10028 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_109
timestamp 1644511149
transform 1 0 11132 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_121
timestamp 1644511149
transform 1 0 12236 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_133
timestamp 1644511149
transform 1 0 13340 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_139
timestamp 1644511149
transform 1 0 13892 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_141
timestamp 1644511149
transform 1 0 14076 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_153
timestamp 1644511149
transform 1 0 15180 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_165
timestamp 1644511149
transform 1 0 16284 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_177
timestamp 1644511149
transform 1 0 17388 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_189
timestamp 1644511149
transform 1 0 18492 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_195
timestamp 1644511149
transform 1 0 19044 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_197
timestamp 1644511149
transform 1 0 19228 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_209
timestamp 1644511149
transform 1 0 20332 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_221
timestamp 1644511149
transform 1 0 21436 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_233
timestamp 1644511149
transform 1 0 22540 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_245
timestamp 1644511149
transform 1 0 23644 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_251
timestamp 1644511149
transform 1 0 24196 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_253
timestamp 1644511149
transform 1 0 24380 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_265
timestamp 1644511149
transform 1 0 25484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_277
timestamp 1644511149
transform 1 0 26588 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_289
timestamp 1644511149
transform 1 0 27692 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_301
timestamp 1644511149
transform 1 0 28796 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_307
timestamp 1644511149
transform 1 0 29348 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_309
timestamp 1644511149
transform 1 0 29532 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_321
timestamp 1644511149
transform 1 0 30636 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_333
timestamp 1644511149
transform 1 0 31740 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_345
timestamp 1644511149
transform 1 0 32844 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_357
timestamp 1644511149
transform 1 0 33948 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_363
timestamp 1644511149
transform 1 0 34500 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_365
timestamp 1644511149
transform 1 0 34684 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_377
timestamp 1644511149
transform 1 0 35788 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_389
timestamp 1644511149
transform 1 0 36892 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_401
timestamp 1644511149
transform 1 0 37996 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_413
timestamp 1644511149
transform 1 0 39100 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_419
timestamp 1644511149
transform 1 0 39652 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_421
timestamp 1644511149
transform 1 0 39836 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_433
timestamp 1644511149
transform 1 0 40940 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_445
timestamp 1644511149
transform 1 0 42044 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_457
timestamp 1644511149
transform 1 0 43148 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_469
timestamp 1644511149
transform 1 0 44252 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_475
timestamp 1644511149
transform 1 0 44804 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_477
timestamp 1644511149
transform 1 0 44988 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_489
timestamp 1644511149
transform 1 0 46092 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_501
timestamp 1644511149
transform 1 0 47196 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_513
timestamp 1644511149
transform 1 0 48300 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_525
timestamp 1644511149
transform 1 0 49404 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_531
timestamp 1644511149
transform 1 0 49956 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_533
timestamp 1644511149
transform 1 0 50140 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_545
timestamp 1644511149
transform 1 0 51244 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_557
timestamp 1644511149
transform 1 0 52348 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_569
timestamp 1644511149
transform 1 0 53452 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_581
timestamp 1644511149
transform 1 0 54556 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_587
timestamp 1644511149
transform 1 0 55108 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_589
timestamp 1644511149
transform 1 0 55292 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_601
timestamp 1644511149
transform 1 0 56396 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_613
timestamp 1644511149
transform 1 0 57500 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_625
timestamp 1644511149
transform 1 0 58604 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_637
timestamp 1644511149
transform 1 0 59708 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_643
timestamp 1644511149
transform 1 0 60260 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_645
timestamp 1644511149
transform 1 0 60444 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_657
timestamp 1644511149
transform 1 0 61548 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_669
timestamp 1644511149
transform 1 0 62652 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_681
timestamp 1644511149
transform 1 0 63756 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_693
timestamp 1644511149
transform 1 0 64860 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_699
timestamp 1644511149
transform 1 0 65412 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_701
timestamp 1644511149
transform 1 0 65596 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_713
timestamp 1644511149
transform 1 0 66700 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_725
timestamp 1644511149
transform 1 0 67804 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_737
timestamp 1644511149
transform 1 0 68908 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_749
timestamp 1644511149
transform 1 0 70012 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_755
timestamp 1644511149
transform 1 0 70564 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_757
timestamp 1644511149
transform 1 0 70748 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_769
timestamp 1644511149
transform 1 0 71852 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_781
timestamp 1644511149
transform 1 0 72956 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_793
timestamp 1644511149
transform 1 0 74060 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_805
timestamp 1644511149
transform 1 0 75164 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_811
timestamp 1644511149
transform 1 0 75716 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_813
timestamp 1644511149
transform 1 0 75900 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_825
timestamp 1644511149
transform 1 0 77004 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_837
timestamp 1644511149
transform 1 0 78108 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_841
timestamp 1644511149
transform 1 0 78476 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_3
timestamp 1644511149
transform 1 0 1380 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_15
timestamp 1644511149
transform 1 0 2484 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_27
timestamp 1644511149
transform 1 0 3588 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_39
timestamp 1644511149
transform 1 0 4692 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_51
timestamp 1644511149
transform 1 0 5796 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_55
timestamp 1644511149
transform 1 0 6164 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_57
timestamp 1644511149
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_69
timestamp 1644511149
transform 1 0 7452 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_81
timestamp 1644511149
transform 1 0 8556 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_93
timestamp 1644511149
transform 1 0 9660 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_105
timestamp 1644511149
transform 1 0 10764 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_111
timestamp 1644511149
transform 1 0 11316 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_113
timestamp 1644511149
transform 1 0 11500 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_125
timestamp 1644511149
transform 1 0 12604 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_137
timestamp 1644511149
transform 1 0 13708 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_149
timestamp 1644511149
transform 1 0 14812 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_161
timestamp 1644511149
transform 1 0 15916 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_167
timestamp 1644511149
transform 1 0 16468 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_169
timestamp 1644511149
transform 1 0 16652 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_181
timestamp 1644511149
transform 1 0 17756 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_193
timestamp 1644511149
transform 1 0 18860 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_205
timestamp 1644511149
transform 1 0 19964 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_217
timestamp 1644511149
transform 1 0 21068 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_223
timestamp 1644511149
transform 1 0 21620 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_225
timestamp 1644511149
transform 1 0 21804 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_237
timestamp 1644511149
transform 1 0 22908 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_249
timestamp 1644511149
transform 1 0 24012 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_261
timestamp 1644511149
transform 1 0 25116 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_273
timestamp 1644511149
transform 1 0 26220 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_279
timestamp 1644511149
transform 1 0 26772 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_281
timestamp 1644511149
transform 1 0 26956 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_293
timestamp 1644511149
transform 1 0 28060 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_305
timestamp 1644511149
transform 1 0 29164 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_317
timestamp 1644511149
transform 1 0 30268 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_329
timestamp 1644511149
transform 1 0 31372 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_335
timestamp 1644511149
transform 1 0 31924 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_337
timestamp 1644511149
transform 1 0 32108 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_349
timestamp 1644511149
transform 1 0 33212 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_361
timestamp 1644511149
transform 1 0 34316 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_373
timestamp 1644511149
transform 1 0 35420 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_385
timestamp 1644511149
transform 1 0 36524 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_391
timestamp 1644511149
transform 1 0 37076 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_393
timestamp 1644511149
transform 1 0 37260 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_405
timestamp 1644511149
transform 1 0 38364 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_417
timestamp 1644511149
transform 1 0 39468 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_429
timestamp 1644511149
transform 1 0 40572 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_441
timestamp 1644511149
transform 1 0 41676 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_447
timestamp 1644511149
transform 1 0 42228 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_449
timestamp 1644511149
transform 1 0 42412 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_461
timestamp 1644511149
transform 1 0 43516 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_473
timestamp 1644511149
transform 1 0 44620 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_485
timestamp 1644511149
transform 1 0 45724 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_497
timestamp 1644511149
transform 1 0 46828 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_503
timestamp 1644511149
transform 1 0 47380 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_505
timestamp 1644511149
transform 1 0 47564 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_517
timestamp 1644511149
transform 1 0 48668 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_529
timestamp 1644511149
transform 1 0 49772 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_541
timestamp 1644511149
transform 1 0 50876 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_553
timestamp 1644511149
transform 1 0 51980 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_559
timestamp 1644511149
transform 1 0 52532 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_561
timestamp 1644511149
transform 1 0 52716 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_573
timestamp 1644511149
transform 1 0 53820 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_585
timestamp 1644511149
transform 1 0 54924 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_597
timestamp 1644511149
transform 1 0 56028 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_609
timestamp 1644511149
transform 1 0 57132 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_615
timestamp 1644511149
transform 1 0 57684 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_617
timestamp 1644511149
transform 1 0 57868 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_629
timestamp 1644511149
transform 1 0 58972 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_641
timestamp 1644511149
transform 1 0 60076 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_653
timestamp 1644511149
transform 1 0 61180 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_665
timestamp 1644511149
transform 1 0 62284 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_671
timestamp 1644511149
transform 1 0 62836 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_673
timestamp 1644511149
transform 1 0 63020 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_685
timestamp 1644511149
transform 1 0 64124 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_697
timestamp 1644511149
transform 1 0 65228 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_709
timestamp 1644511149
transform 1 0 66332 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_721
timestamp 1644511149
transform 1 0 67436 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_727
timestamp 1644511149
transform 1 0 67988 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_729
timestamp 1644511149
transform 1 0 68172 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_741
timestamp 1644511149
transform 1 0 69276 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_753
timestamp 1644511149
transform 1 0 70380 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_765
timestamp 1644511149
transform 1 0 71484 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_777
timestamp 1644511149
transform 1 0 72588 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_783
timestamp 1644511149
transform 1 0 73140 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_785
timestamp 1644511149
transform 1 0 73324 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_797
timestamp 1644511149
transform 1 0 74428 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_809
timestamp 1644511149
transform 1 0 75532 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_821
timestamp 1644511149
transform 1 0 76636 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_833
timestamp 1644511149
transform 1 0 77740 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_839
timestamp 1644511149
transform 1 0 78292 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_53_841
timestamp 1644511149
transform 1 0 78476 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_9
timestamp 1644511149
transform 1 0 1932 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_21
timestamp 1644511149
transform 1 0 3036 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_27
timestamp 1644511149
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_29
timestamp 1644511149
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_41
timestamp 1644511149
transform 1 0 4876 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_53
timestamp 1644511149
transform 1 0 5980 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_65
timestamp 1644511149
transform 1 0 7084 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_77
timestamp 1644511149
transform 1 0 8188 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_83
timestamp 1644511149
transform 1 0 8740 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_85
timestamp 1644511149
transform 1 0 8924 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_97
timestamp 1644511149
transform 1 0 10028 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_109
timestamp 1644511149
transform 1 0 11132 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_121
timestamp 1644511149
transform 1 0 12236 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_133
timestamp 1644511149
transform 1 0 13340 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_139
timestamp 1644511149
transform 1 0 13892 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_141
timestamp 1644511149
transform 1 0 14076 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_153
timestamp 1644511149
transform 1 0 15180 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_165
timestamp 1644511149
transform 1 0 16284 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_177
timestamp 1644511149
transform 1 0 17388 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_189
timestamp 1644511149
transform 1 0 18492 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_195
timestamp 1644511149
transform 1 0 19044 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_197
timestamp 1644511149
transform 1 0 19228 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_209
timestamp 1644511149
transform 1 0 20332 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_221
timestamp 1644511149
transform 1 0 21436 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_233
timestamp 1644511149
transform 1 0 22540 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_245
timestamp 1644511149
transform 1 0 23644 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_251
timestamp 1644511149
transform 1 0 24196 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_253
timestamp 1644511149
transform 1 0 24380 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_265
timestamp 1644511149
transform 1 0 25484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_277
timestamp 1644511149
transform 1 0 26588 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_289
timestamp 1644511149
transform 1 0 27692 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_301
timestamp 1644511149
transform 1 0 28796 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_307
timestamp 1644511149
transform 1 0 29348 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_309
timestamp 1644511149
transform 1 0 29532 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_321
timestamp 1644511149
transform 1 0 30636 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_333
timestamp 1644511149
transform 1 0 31740 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_345
timestamp 1644511149
transform 1 0 32844 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_357
timestamp 1644511149
transform 1 0 33948 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_363
timestamp 1644511149
transform 1 0 34500 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_365
timestamp 1644511149
transform 1 0 34684 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_377
timestamp 1644511149
transform 1 0 35788 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_389
timestamp 1644511149
transform 1 0 36892 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_401
timestamp 1644511149
transform 1 0 37996 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_413
timestamp 1644511149
transform 1 0 39100 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_419
timestamp 1644511149
transform 1 0 39652 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_421
timestamp 1644511149
transform 1 0 39836 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_433
timestamp 1644511149
transform 1 0 40940 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_445
timestamp 1644511149
transform 1 0 42044 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_457
timestamp 1644511149
transform 1 0 43148 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_469
timestamp 1644511149
transform 1 0 44252 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_475
timestamp 1644511149
transform 1 0 44804 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_477
timestamp 1644511149
transform 1 0 44988 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_489
timestamp 1644511149
transform 1 0 46092 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_501
timestamp 1644511149
transform 1 0 47196 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_513
timestamp 1644511149
transform 1 0 48300 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_525
timestamp 1644511149
transform 1 0 49404 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_531
timestamp 1644511149
transform 1 0 49956 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_533
timestamp 1644511149
transform 1 0 50140 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_545
timestamp 1644511149
transform 1 0 51244 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_557
timestamp 1644511149
transform 1 0 52348 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_569
timestamp 1644511149
transform 1 0 53452 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_581
timestamp 1644511149
transform 1 0 54556 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_587
timestamp 1644511149
transform 1 0 55108 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_589
timestamp 1644511149
transform 1 0 55292 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_601
timestamp 1644511149
transform 1 0 56396 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_613
timestamp 1644511149
transform 1 0 57500 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_625
timestamp 1644511149
transform 1 0 58604 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_637
timestamp 1644511149
transform 1 0 59708 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_643
timestamp 1644511149
transform 1 0 60260 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_645
timestamp 1644511149
transform 1 0 60444 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_657
timestamp 1644511149
transform 1 0 61548 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_669
timestamp 1644511149
transform 1 0 62652 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_681
timestamp 1644511149
transform 1 0 63756 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_693
timestamp 1644511149
transform 1 0 64860 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_699
timestamp 1644511149
transform 1 0 65412 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_701
timestamp 1644511149
transform 1 0 65596 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_713
timestamp 1644511149
transform 1 0 66700 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_725
timestamp 1644511149
transform 1 0 67804 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_737
timestamp 1644511149
transform 1 0 68908 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_749
timestamp 1644511149
transform 1 0 70012 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_755
timestamp 1644511149
transform 1 0 70564 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_757
timestamp 1644511149
transform 1 0 70748 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_769
timestamp 1644511149
transform 1 0 71852 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_781
timestamp 1644511149
transform 1 0 72956 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_793
timestamp 1644511149
transform 1 0 74060 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_805
timestamp 1644511149
transform 1 0 75164 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_811
timestamp 1644511149
transform 1 0 75716 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_813
timestamp 1644511149
transform 1 0 75900 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_825
timestamp 1644511149
transform 1 0 77004 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_54_837
timestamp 1644511149
transform 1 0 78108 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_841
timestamp 1644511149
transform 1 0 78476 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_3
timestamp 1644511149
transform 1 0 1380 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_15
timestamp 1644511149
transform 1 0 2484 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_27
timestamp 1644511149
transform 1 0 3588 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_39
timestamp 1644511149
transform 1 0 4692 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_51
timestamp 1644511149
transform 1 0 5796 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_55
timestamp 1644511149
transform 1 0 6164 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_57
timestamp 1644511149
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_69
timestamp 1644511149
transform 1 0 7452 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_81
timestamp 1644511149
transform 1 0 8556 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_93
timestamp 1644511149
transform 1 0 9660 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_105
timestamp 1644511149
transform 1 0 10764 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_111
timestamp 1644511149
transform 1 0 11316 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_113
timestamp 1644511149
transform 1 0 11500 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_125
timestamp 1644511149
transform 1 0 12604 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_137
timestamp 1644511149
transform 1 0 13708 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_149
timestamp 1644511149
transform 1 0 14812 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_161
timestamp 1644511149
transform 1 0 15916 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_167
timestamp 1644511149
transform 1 0 16468 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_169
timestamp 1644511149
transform 1 0 16652 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_181
timestamp 1644511149
transform 1 0 17756 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_193
timestamp 1644511149
transform 1 0 18860 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_205
timestamp 1644511149
transform 1 0 19964 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_217
timestamp 1644511149
transform 1 0 21068 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_223
timestamp 1644511149
transform 1 0 21620 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_225
timestamp 1644511149
transform 1 0 21804 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_237
timestamp 1644511149
transform 1 0 22908 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_249
timestamp 1644511149
transform 1 0 24012 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_261
timestamp 1644511149
transform 1 0 25116 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_273
timestamp 1644511149
transform 1 0 26220 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_279
timestamp 1644511149
transform 1 0 26772 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_281
timestamp 1644511149
transform 1 0 26956 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_293
timestamp 1644511149
transform 1 0 28060 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_305
timestamp 1644511149
transform 1 0 29164 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_317
timestamp 1644511149
transform 1 0 30268 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_329
timestamp 1644511149
transform 1 0 31372 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_335
timestamp 1644511149
transform 1 0 31924 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_337
timestamp 1644511149
transform 1 0 32108 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_349
timestamp 1644511149
transform 1 0 33212 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_361
timestamp 1644511149
transform 1 0 34316 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_373
timestamp 1644511149
transform 1 0 35420 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_385
timestamp 1644511149
transform 1 0 36524 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_391
timestamp 1644511149
transform 1 0 37076 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_393
timestamp 1644511149
transform 1 0 37260 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_405
timestamp 1644511149
transform 1 0 38364 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_417
timestamp 1644511149
transform 1 0 39468 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_429
timestamp 1644511149
transform 1 0 40572 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_441
timestamp 1644511149
transform 1 0 41676 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_447
timestamp 1644511149
transform 1 0 42228 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_449
timestamp 1644511149
transform 1 0 42412 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_461
timestamp 1644511149
transform 1 0 43516 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_473
timestamp 1644511149
transform 1 0 44620 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_485
timestamp 1644511149
transform 1 0 45724 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_497
timestamp 1644511149
transform 1 0 46828 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_503
timestamp 1644511149
transform 1 0 47380 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_505
timestamp 1644511149
transform 1 0 47564 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_517
timestamp 1644511149
transform 1 0 48668 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_529
timestamp 1644511149
transform 1 0 49772 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_541
timestamp 1644511149
transform 1 0 50876 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_553
timestamp 1644511149
transform 1 0 51980 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_559
timestamp 1644511149
transform 1 0 52532 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_561
timestamp 1644511149
transform 1 0 52716 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_573
timestamp 1644511149
transform 1 0 53820 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_585
timestamp 1644511149
transform 1 0 54924 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_597
timestamp 1644511149
transform 1 0 56028 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_609
timestamp 1644511149
transform 1 0 57132 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_615
timestamp 1644511149
transform 1 0 57684 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_617
timestamp 1644511149
transform 1 0 57868 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_629
timestamp 1644511149
transform 1 0 58972 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_641
timestamp 1644511149
transform 1 0 60076 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_653
timestamp 1644511149
transform 1 0 61180 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_665
timestamp 1644511149
transform 1 0 62284 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_671
timestamp 1644511149
transform 1 0 62836 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_673
timestamp 1644511149
transform 1 0 63020 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_685
timestamp 1644511149
transform 1 0 64124 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_697
timestamp 1644511149
transform 1 0 65228 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_709
timestamp 1644511149
transform 1 0 66332 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_721
timestamp 1644511149
transform 1 0 67436 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_727
timestamp 1644511149
transform 1 0 67988 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_729
timestamp 1644511149
transform 1 0 68172 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_741
timestamp 1644511149
transform 1 0 69276 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_753
timestamp 1644511149
transform 1 0 70380 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_765
timestamp 1644511149
transform 1 0 71484 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_777
timestamp 1644511149
transform 1 0 72588 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_783
timestamp 1644511149
transform 1 0 73140 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_785
timestamp 1644511149
transform 1 0 73324 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_797
timestamp 1644511149
transform 1 0 74428 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_809
timestamp 1644511149
transform 1 0 75532 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_821
timestamp 1644511149
transform 1 0 76636 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_55_829
timestamp 1644511149
transform 1 0 77372 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_55_836
timestamp 1644511149
transform 1 0 78016 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_841
timestamp 1644511149
transform 1 0 78476 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_3
timestamp 1644511149
transform 1 0 1380 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_15
timestamp 1644511149
transform 1 0 2484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_27
timestamp 1644511149
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_29
timestamp 1644511149
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_41
timestamp 1644511149
transform 1 0 4876 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_53
timestamp 1644511149
transform 1 0 5980 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_65
timestamp 1644511149
transform 1 0 7084 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_77
timestamp 1644511149
transform 1 0 8188 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_83
timestamp 1644511149
transform 1 0 8740 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_85
timestamp 1644511149
transform 1 0 8924 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_97
timestamp 1644511149
transform 1 0 10028 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_109
timestamp 1644511149
transform 1 0 11132 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_121
timestamp 1644511149
transform 1 0 12236 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_133
timestamp 1644511149
transform 1 0 13340 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_139
timestamp 1644511149
transform 1 0 13892 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_141
timestamp 1644511149
transform 1 0 14076 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_153
timestamp 1644511149
transform 1 0 15180 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_165
timestamp 1644511149
transform 1 0 16284 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_177
timestamp 1644511149
transform 1 0 17388 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_189
timestamp 1644511149
transform 1 0 18492 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_195
timestamp 1644511149
transform 1 0 19044 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_197
timestamp 1644511149
transform 1 0 19228 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_209
timestamp 1644511149
transform 1 0 20332 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_221
timestamp 1644511149
transform 1 0 21436 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_233
timestamp 1644511149
transform 1 0 22540 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_245
timestamp 1644511149
transform 1 0 23644 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_251
timestamp 1644511149
transform 1 0 24196 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_253
timestamp 1644511149
transform 1 0 24380 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_265
timestamp 1644511149
transform 1 0 25484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_277
timestamp 1644511149
transform 1 0 26588 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_289
timestamp 1644511149
transform 1 0 27692 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_301
timestamp 1644511149
transform 1 0 28796 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_307
timestamp 1644511149
transform 1 0 29348 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_309
timestamp 1644511149
transform 1 0 29532 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_321
timestamp 1644511149
transform 1 0 30636 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_333
timestamp 1644511149
transform 1 0 31740 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_345
timestamp 1644511149
transform 1 0 32844 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_357
timestamp 1644511149
transform 1 0 33948 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_363
timestamp 1644511149
transform 1 0 34500 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_365
timestamp 1644511149
transform 1 0 34684 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_377
timestamp 1644511149
transform 1 0 35788 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_389
timestamp 1644511149
transform 1 0 36892 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_401
timestamp 1644511149
transform 1 0 37996 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_413
timestamp 1644511149
transform 1 0 39100 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_419
timestamp 1644511149
transform 1 0 39652 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_421
timestamp 1644511149
transform 1 0 39836 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_433
timestamp 1644511149
transform 1 0 40940 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_445
timestamp 1644511149
transform 1 0 42044 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_457
timestamp 1644511149
transform 1 0 43148 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_469
timestamp 1644511149
transform 1 0 44252 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_475
timestamp 1644511149
transform 1 0 44804 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_477
timestamp 1644511149
transform 1 0 44988 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_489
timestamp 1644511149
transform 1 0 46092 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_501
timestamp 1644511149
transform 1 0 47196 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_513
timestamp 1644511149
transform 1 0 48300 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_525
timestamp 1644511149
transform 1 0 49404 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_531
timestamp 1644511149
transform 1 0 49956 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_533
timestamp 1644511149
transform 1 0 50140 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_545
timestamp 1644511149
transform 1 0 51244 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_557
timestamp 1644511149
transform 1 0 52348 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_569
timestamp 1644511149
transform 1 0 53452 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_581
timestamp 1644511149
transform 1 0 54556 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_587
timestamp 1644511149
transform 1 0 55108 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_589
timestamp 1644511149
transform 1 0 55292 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_601
timestamp 1644511149
transform 1 0 56396 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_613
timestamp 1644511149
transform 1 0 57500 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_625
timestamp 1644511149
transform 1 0 58604 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_637
timestamp 1644511149
transform 1 0 59708 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_643
timestamp 1644511149
transform 1 0 60260 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_645
timestamp 1644511149
transform 1 0 60444 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_657
timestamp 1644511149
transform 1 0 61548 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_669
timestamp 1644511149
transform 1 0 62652 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_681
timestamp 1644511149
transform 1 0 63756 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_693
timestamp 1644511149
transform 1 0 64860 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_699
timestamp 1644511149
transform 1 0 65412 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_701
timestamp 1644511149
transform 1 0 65596 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_713
timestamp 1644511149
transform 1 0 66700 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_725
timestamp 1644511149
transform 1 0 67804 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_737
timestamp 1644511149
transform 1 0 68908 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_749
timestamp 1644511149
transform 1 0 70012 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_755
timestamp 1644511149
transform 1 0 70564 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_757
timestamp 1644511149
transform 1 0 70748 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_769
timestamp 1644511149
transform 1 0 71852 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_781
timestamp 1644511149
transform 1 0 72956 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_793
timestamp 1644511149
transform 1 0 74060 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_805
timestamp 1644511149
transform 1 0 75164 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_811
timestamp 1644511149
transform 1 0 75716 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_813
timestamp 1644511149
transform 1 0 75900 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_825
timestamp 1644511149
transform 1 0 77004 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_56_833
timestamp 1644511149
transform 1 0 77740 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_837
timestamp 1644511149
transform 1 0 78108 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_841
timestamp 1644511149
transform 1 0 78476 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_3
timestamp 1644511149
transform 1 0 1380 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_15
timestamp 1644511149
transform 1 0 2484 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_27
timestamp 1644511149
transform 1 0 3588 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_39
timestamp 1644511149
transform 1 0 4692 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_51
timestamp 1644511149
transform 1 0 5796 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_55
timestamp 1644511149
transform 1 0 6164 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_57
timestamp 1644511149
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_69
timestamp 1644511149
transform 1 0 7452 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_81
timestamp 1644511149
transform 1 0 8556 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_93
timestamp 1644511149
transform 1 0 9660 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_105
timestamp 1644511149
transform 1 0 10764 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_111
timestamp 1644511149
transform 1 0 11316 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_113
timestamp 1644511149
transform 1 0 11500 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_125
timestamp 1644511149
transform 1 0 12604 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_137
timestamp 1644511149
transform 1 0 13708 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_149
timestamp 1644511149
transform 1 0 14812 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_161
timestamp 1644511149
transform 1 0 15916 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_167
timestamp 1644511149
transform 1 0 16468 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_169
timestamp 1644511149
transform 1 0 16652 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_181
timestamp 1644511149
transform 1 0 17756 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_193
timestamp 1644511149
transform 1 0 18860 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_205
timestamp 1644511149
transform 1 0 19964 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_217
timestamp 1644511149
transform 1 0 21068 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_223
timestamp 1644511149
transform 1 0 21620 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_225
timestamp 1644511149
transform 1 0 21804 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_237
timestamp 1644511149
transform 1 0 22908 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_249
timestamp 1644511149
transform 1 0 24012 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_261
timestamp 1644511149
transform 1 0 25116 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_273
timestamp 1644511149
transform 1 0 26220 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_279
timestamp 1644511149
transform 1 0 26772 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_281
timestamp 1644511149
transform 1 0 26956 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_293
timestamp 1644511149
transform 1 0 28060 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_305
timestamp 1644511149
transform 1 0 29164 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_317
timestamp 1644511149
transform 1 0 30268 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_329
timestamp 1644511149
transform 1 0 31372 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_335
timestamp 1644511149
transform 1 0 31924 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_337
timestamp 1644511149
transform 1 0 32108 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_349
timestamp 1644511149
transform 1 0 33212 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_361
timestamp 1644511149
transform 1 0 34316 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_373
timestamp 1644511149
transform 1 0 35420 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_385
timestamp 1644511149
transform 1 0 36524 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_391
timestamp 1644511149
transform 1 0 37076 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_393
timestamp 1644511149
transform 1 0 37260 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_405
timestamp 1644511149
transform 1 0 38364 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_417
timestamp 1644511149
transform 1 0 39468 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_429
timestamp 1644511149
transform 1 0 40572 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_441
timestamp 1644511149
transform 1 0 41676 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_447
timestamp 1644511149
transform 1 0 42228 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_449
timestamp 1644511149
transform 1 0 42412 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_461
timestamp 1644511149
transform 1 0 43516 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_473
timestamp 1644511149
transform 1 0 44620 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_485
timestamp 1644511149
transform 1 0 45724 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_497
timestamp 1644511149
transform 1 0 46828 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_503
timestamp 1644511149
transform 1 0 47380 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_505
timestamp 1644511149
transform 1 0 47564 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_517
timestamp 1644511149
transform 1 0 48668 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_529
timestamp 1644511149
transform 1 0 49772 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_541
timestamp 1644511149
transform 1 0 50876 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_553
timestamp 1644511149
transform 1 0 51980 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_559
timestamp 1644511149
transform 1 0 52532 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_561
timestamp 1644511149
transform 1 0 52716 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_573
timestamp 1644511149
transform 1 0 53820 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_585
timestamp 1644511149
transform 1 0 54924 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_597
timestamp 1644511149
transform 1 0 56028 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_609
timestamp 1644511149
transform 1 0 57132 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_615
timestamp 1644511149
transform 1 0 57684 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_617
timestamp 1644511149
transform 1 0 57868 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_629
timestamp 1644511149
transform 1 0 58972 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_641
timestamp 1644511149
transform 1 0 60076 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_653
timestamp 1644511149
transform 1 0 61180 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_665
timestamp 1644511149
transform 1 0 62284 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_671
timestamp 1644511149
transform 1 0 62836 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_673
timestamp 1644511149
transform 1 0 63020 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_685
timestamp 1644511149
transform 1 0 64124 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_697
timestamp 1644511149
transform 1 0 65228 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_709
timestamp 1644511149
transform 1 0 66332 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_721
timestamp 1644511149
transform 1 0 67436 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_727
timestamp 1644511149
transform 1 0 67988 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_729
timestamp 1644511149
transform 1 0 68172 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_741
timestamp 1644511149
transform 1 0 69276 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_753
timestamp 1644511149
transform 1 0 70380 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_765
timestamp 1644511149
transform 1 0 71484 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_777
timestamp 1644511149
transform 1 0 72588 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_783
timestamp 1644511149
transform 1 0 73140 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_785
timestamp 1644511149
transform 1 0 73324 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_797
timestamp 1644511149
transform 1 0 74428 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_809
timestamp 1644511149
transform 1 0 75532 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_821
timestamp 1644511149
transform 1 0 76636 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_833
timestamp 1644511149
transform 1 0 77740 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_839
timestamp 1644511149
transform 1 0 78292 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_57_841
timestamp 1644511149
transform 1 0 78476 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_3
timestamp 1644511149
transform 1 0 1380 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_15
timestamp 1644511149
transform 1 0 2484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_27
timestamp 1644511149
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_29
timestamp 1644511149
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_41
timestamp 1644511149
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_53
timestamp 1644511149
transform 1 0 5980 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_65
timestamp 1644511149
transform 1 0 7084 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_77
timestamp 1644511149
transform 1 0 8188 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_83
timestamp 1644511149
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_85
timestamp 1644511149
transform 1 0 8924 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_97
timestamp 1644511149
transform 1 0 10028 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_109
timestamp 1644511149
transform 1 0 11132 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_121
timestamp 1644511149
transform 1 0 12236 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_133
timestamp 1644511149
transform 1 0 13340 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_139
timestamp 1644511149
transform 1 0 13892 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_141
timestamp 1644511149
transform 1 0 14076 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_153
timestamp 1644511149
transform 1 0 15180 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_165
timestamp 1644511149
transform 1 0 16284 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_177
timestamp 1644511149
transform 1 0 17388 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_189
timestamp 1644511149
transform 1 0 18492 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_195
timestamp 1644511149
transform 1 0 19044 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_197
timestamp 1644511149
transform 1 0 19228 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_209
timestamp 1644511149
transform 1 0 20332 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_221
timestamp 1644511149
transform 1 0 21436 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_233
timestamp 1644511149
transform 1 0 22540 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_245
timestamp 1644511149
transform 1 0 23644 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_251
timestamp 1644511149
transform 1 0 24196 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_253
timestamp 1644511149
transform 1 0 24380 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_265
timestamp 1644511149
transform 1 0 25484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_277
timestamp 1644511149
transform 1 0 26588 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_289
timestamp 1644511149
transform 1 0 27692 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_301
timestamp 1644511149
transform 1 0 28796 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_307
timestamp 1644511149
transform 1 0 29348 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_309
timestamp 1644511149
transform 1 0 29532 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_321
timestamp 1644511149
transform 1 0 30636 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_333
timestamp 1644511149
transform 1 0 31740 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_345
timestamp 1644511149
transform 1 0 32844 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_357
timestamp 1644511149
transform 1 0 33948 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_363
timestamp 1644511149
transform 1 0 34500 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_365
timestamp 1644511149
transform 1 0 34684 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_377
timestamp 1644511149
transform 1 0 35788 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_389
timestamp 1644511149
transform 1 0 36892 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_401
timestamp 1644511149
transform 1 0 37996 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_413
timestamp 1644511149
transform 1 0 39100 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_419
timestamp 1644511149
transform 1 0 39652 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_421
timestamp 1644511149
transform 1 0 39836 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_433
timestamp 1644511149
transform 1 0 40940 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_445
timestamp 1644511149
transform 1 0 42044 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_457
timestamp 1644511149
transform 1 0 43148 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_469
timestamp 1644511149
transform 1 0 44252 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_475
timestamp 1644511149
transform 1 0 44804 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_477
timestamp 1644511149
transform 1 0 44988 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_489
timestamp 1644511149
transform 1 0 46092 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_501
timestamp 1644511149
transform 1 0 47196 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_513
timestamp 1644511149
transform 1 0 48300 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_525
timestamp 1644511149
transform 1 0 49404 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_531
timestamp 1644511149
transform 1 0 49956 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_533
timestamp 1644511149
transform 1 0 50140 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_545
timestamp 1644511149
transform 1 0 51244 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_557
timestamp 1644511149
transform 1 0 52348 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_569
timestamp 1644511149
transform 1 0 53452 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_581
timestamp 1644511149
transform 1 0 54556 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_587
timestamp 1644511149
transform 1 0 55108 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_589
timestamp 1644511149
transform 1 0 55292 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_601
timestamp 1644511149
transform 1 0 56396 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_613
timestamp 1644511149
transform 1 0 57500 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_625
timestamp 1644511149
transform 1 0 58604 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_637
timestamp 1644511149
transform 1 0 59708 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_643
timestamp 1644511149
transform 1 0 60260 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_645
timestamp 1644511149
transform 1 0 60444 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_657
timestamp 1644511149
transform 1 0 61548 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_669
timestamp 1644511149
transform 1 0 62652 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_681
timestamp 1644511149
transform 1 0 63756 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_693
timestamp 1644511149
transform 1 0 64860 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_699
timestamp 1644511149
transform 1 0 65412 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_701
timestamp 1644511149
transform 1 0 65596 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_713
timestamp 1644511149
transform 1 0 66700 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_725
timestamp 1644511149
transform 1 0 67804 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_737
timestamp 1644511149
transform 1 0 68908 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_749
timestamp 1644511149
transform 1 0 70012 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_755
timestamp 1644511149
transform 1 0 70564 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_757
timestamp 1644511149
transform 1 0 70748 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_769
timestamp 1644511149
transform 1 0 71852 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_781
timestamp 1644511149
transform 1 0 72956 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_793
timestamp 1644511149
transform 1 0 74060 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_805
timestamp 1644511149
transform 1 0 75164 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_811
timestamp 1644511149
transform 1 0 75716 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_813
timestamp 1644511149
transform 1 0 75900 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_825
timestamp 1644511149
transform 1 0 77004 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_58_837
timestamp 1644511149
transform 1 0 78108 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_841
timestamp 1644511149
transform 1 0 78476 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_3
timestamp 1644511149
transform 1 0 1380 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_15
timestamp 1644511149
transform 1 0 2484 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_27
timestamp 1644511149
transform 1 0 3588 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_39
timestamp 1644511149
transform 1 0 4692 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_51
timestamp 1644511149
transform 1 0 5796 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_55
timestamp 1644511149
transform 1 0 6164 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_57
timestamp 1644511149
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_69
timestamp 1644511149
transform 1 0 7452 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_81
timestamp 1644511149
transform 1 0 8556 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_93
timestamp 1644511149
transform 1 0 9660 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_105
timestamp 1644511149
transform 1 0 10764 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_111
timestamp 1644511149
transform 1 0 11316 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_113
timestamp 1644511149
transform 1 0 11500 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_125
timestamp 1644511149
transform 1 0 12604 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_137
timestamp 1644511149
transform 1 0 13708 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_149
timestamp 1644511149
transform 1 0 14812 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_161
timestamp 1644511149
transform 1 0 15916 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_167
timestamp 1644511149
transform 1 0 16468 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_169
timestamp 1644511149
transform 1 0 16652 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_181
timestamp 1644511149
transform 1 0 17756 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_193
timestamp 1644511149
transform 1 0 18860 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_205
timestamp 1644511149
transform 1 0 19964 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_217
timestamp 1644511149
transform 1 0 21068 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_223
timestamp 1644511149
transform 1 0 21620 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_225
timestamp 1644511149
transform 1 0 21804 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_237
timestamp 1644511149
transform 1 0 22908 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_249
timestamp 1644511149
transform 1 0 24012 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_261
timestamp 1644511149
transform 1 0 25116 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_273
timestamp 1644511149
transform 1 0 26220 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_279
timestamp 1644511149
transform 1 0 26772 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_281
timestamp 1644511149
transform 1 0 26956 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_293
timestamp 1644511149
transform 1 0 28060 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_305
timestamp 1644511149
transform 1 0 29164 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_317
timestamp 1644511149
transform 1 0 30268 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_329
timestamp 1644511149
transform 1 0 31372 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_335
timestamp 1644511149
transform 1 0 31924 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_337
timestamp 1644511149
transform 1 0 32108 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_349
timestamp 1644511149
transform 1 0 33212 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_361
timestamp 1644511149
transform 1 0 34316 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_373
timestamp 1644511149
transform 1 0 35420 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_385
timestamp 1644511149
transform 1 0 36524 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_391
timestamp 1644511149
transform 1 0 37076 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_393
timestamp 1644511149
transform 1 0 37260 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_405
timestamp 1644511149
transform 1 0 38364 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_417
timestamp 1644511149
transform 1 0 39468 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_429
timestamp 1644511149
transform 1 0 40572 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_441
timestamp 1644511149
transform 1 0 41676 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_447
timestamp 1644511149
transform 1 0 42228 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_449
timestamp 1644511149
transform 1 0 42412 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_461
timestamp 1644511149
transform 1 0 43516 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_473
timestamp 1644511149
transform 1 0 44620 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_485
timestamp 1644511149
transform 1 0 45724 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_497
timestamp 1644511149
transform 1 0 46828 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_503
timestamp 1644511149
transform 1 0 47380 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_505
timestamp 1644511149
transform 1 0 47564 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_517
timestamp 1644511149
transform 1 0 48668 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_529
timestamp 1644511149
transform 1 0 49772 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_541
timestamp 1644511149
transform 1 0 50876 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_553
timestamp 1644511149
transform 1 0 51980 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_559
timestamp 1644511149
transform 1 0 52532 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_561
timestamp 1644511149
transform 1 0 52716 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_573
timestamp 1644511149
transform 1 0 53820 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_585
timestamp 1644511149
transform 1 0 54924 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_597
timestamp 1644511149
transform 1 0 56028 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_609
timestamp 1644511149
transform 1 0 57132 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_615
timestamp 1644511149
transform 1 0 57684 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_617
timestamp 1644511149
transform 1 0 57868 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_629
timestamp 1644511149
transform 1 0 58972 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_641
timestamp 1644511149
transform 1 0 60076 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_653
timestamp 1644511149
transform 1 0 61180 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_665
timestamp 1644511149
transform 1 0 62284 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_671
timestamp 1644511149
transform 1 0 62836 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_673
timestamp 1644511149
transform 1 0 63020 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_685
timestamp 1644511149
transform 1 0 64124 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_697
timestamp 1644511149
transform 1 0 65228 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_709
timestamp 1644511149
transform 1 0 66332 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_721
timestamp 1644511149
transform 1 0 67436 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_727
timestamp 1644511149
transform 1 0 67988 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_729
timestamp 1644511149
transform 1 0 68172 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_741
timestamp 1644511149
transform 1 0 69276 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_753
timestamp 1644511149
transform 1 0 70380 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_59_765
timestamp 1644511149
transform 1 0 71484 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_770
timestamp 1644511149
transform 1 0 71944 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_59_782
timestamp 1644511149
transform 1 0 73048 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_59_785
timestamp 1644511149
transform 1 0 73324 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_797
timestamp 1644511149
transform 1 0 74428 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_809
timestamp 1644511149
transform 1 0 75532 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_821
timestamp 1644511149
transform 1 0 76636 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_833
timestamp 1644511149
transform 1 0 77740 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_839
timestamp 1644511149
transform 1 0 78292 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_59_841
timestamp 1644511149
transform 1 0 78476 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_7
timestamp 1644511149
transform 1 0 1748 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_19
timestamp 1644511149
transform 1 0 2852 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_60_27
timestamp 1644511149
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_29
timestamp 1644511149
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_41
timestamp 1644511149
transform 1 0 4876 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_53
timestamp 1644511149
transform 1 0 5980 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_65
timestamp 1644511149
transform 1 0 7084 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_77
timestamp 1644511149
transform 1 0 8188 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_83
timestamp 1644511149
transform 1 0 8740 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_85
timestamp 1644511149
transform 1 0 8924 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_97
timestamp 1644511149
transform 1 0 10028 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_109
timestamp 1644511149
transform 1 0 11132 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_121
timestamp 1644511149
transform 1 0 12236 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_133
timestamp 1644511149
transform 1 0 13340 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_139
timestamp 1644511149
transform 1 0 13892 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_141
timestamp 1644511149
transform 1 0 14076 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_153
timestamp 1644511149
transform 1 0 15180 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_165
timestamp 1644511149
transform 1 0 16284 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_177
timestamp 1644511149
transform 1 0 17388 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_189
timestamp 1644511149
transform 1 0 18492 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_195
timestamp 1644511149
transform 1 0 19044 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_197
timestamp 1644511149
transform 1 0 19228 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_209
timestamp 1644511149
transform 1 0 20332 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_221
timestamp 1644511149
transform 1 0 21436 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_233
timestamp 1644511149
transform 1 0 22540 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_245
timestamp 1644511149
transform 1 0 23644 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_251
timestamp 1644511149
transform 1 0 24196 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_253
timestamp 1644511149
transform 1 0 24380 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_265
timestamp 1644511149
transform 1 0 25484 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_277
timestamp 1644511149
transform 1 0 26588 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_289
timestamp 1644511149
transform 1 0 27692 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_301
timestamp 1644511149
transform 1 0 28796 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_307
timestamp 1644511149
transform 1 0 29348 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_309
timestamp 1644511149
transform 1 0 29532 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_321
timestamp 1644511149
transform 1 0 30636 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_333
timestamp 1644511149
transform 1 0 31740 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_345
timestamp 1644511149
transform 1 0 32844 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_357
timestamp 1644511149
transform 1 0 33948 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_363
timestamp 1644511149
transform 1 0 34500 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_365
timestamp 1644511149
transform 1 0 34684 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_377
timestamp 1644511149
transform 1 0 35788 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_389
timestamp 1644511149
transform 1 0 36892 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_401
timestamp 1644511149
transform 1 0 37996 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_413
timestamp 1644511149
transform 1 0 39100 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_419
timestamp 1644511149
transform 1 0 39652 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_421
timestamp 1644511149
transform 1 0 39836 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_433
timestamp 1644511149
transform 1 0 40940 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_445
timestamp 1644511149
transform 1 0 42044 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_457
timestamp 1644511149
transform 1 0 43148 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_469
timestamp 1644511149
transform 1 0 44252 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_475
timestamp 1644511149
transform 1 0 44804 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_477
timestamp 1644511149
transform 1 0 44988 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_489
timestamp 1644511149
transform 1 0 46092 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_501
timestamp 1644511149
transform 1 0 47196 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_513
timestamp 1644511149
transform 1 0 48300 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_525
timestamp 1644511149
transform 1 0 49404 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_531
timestamp 1644511149
transform 1 0 49956 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_533
timestamp 1644511149
transform 1 0 50140 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_545
timestamp 1644511149
transform 1 0 51244 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_557
timestamp 1644511149
transform 1 0 52348 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_569
timestamp 1644511149
transform 1 0 53452 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_581
timestamp 1644511149
transform 1 0 54556 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_587
timestamp 1644511149
transform 1 0 55108 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_589
timestamp 1644511149
transform 1 0 55292 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_601
timestamp 1644511149
transform 1 0 56396 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_613
timestamp 1644511149
transform 1 0 57500 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_625
timestamp 1644511149
transform 1 0 58604 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_637
timestamp 1644511149
transform 1 0 59708 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_643
timestamp 1644511149
transform 1 0 60260 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_645
timestamp 1644511149
transform 1 0 60444 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_657
timestamp 1644511149
transform 1 0 61548 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_669
timestamp 1644511149
transform 1 0 62652 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_681
timestamp 1644511149
transform 1 0 63756 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_693
timestamp 1644511149
transform 1 0 64860 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_699
timestamp 1644511149
transform 1 0 65412 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_701
timestamp 1644511149
transform 1 0 65596 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_713
timestamp 1644511149
transform 1 0 66700 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_725
timestamp 1644511149
transform 1 0 67804 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_737
timestamp 1644511149
transform 1 0 68908 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_749
timestamp 1644511149
transform 1 0 70012 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_755
timestamp 1644511149
transform 1 0 70564 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_757
timestamp 1644511149
transform 1 0 70748 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_769
timestamp 1644511149
transform 1 0 71852 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_781
timestamp 1644511149
transform 1 0 72956 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_793
timestamp 1644511149
transform 1 0 74060 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_805
timestamp 1644511149
transform 1 0 75164 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_811
timestamp 1644511149
transform 1 0 75716 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_813
timestamp 1644511149
transform 1 0 75900 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_825
timestamp 1644511149
transform 1 0 77004 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_837
timestamp 1644511149
transform 1 0 78108 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_841
timestamp 1644511149
transform 1 0 78476 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_3
timestamp 1644511149
transform 1 0 1380 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_15
timestamp 1644511149
transform 1 0 2484 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_27
timestamp 1644511149
transform 1 0 3588 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_39
timestamp 1644511149
transform 1 0 4692 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_51
timestamp 1644511149
transform 1 0 5796 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_55
timestamp 1644511149
transform 1 0 6164 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_57
timestamp 1644511149
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_69
timestamp 1644511149
transform 1 0 7452 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_81
timestamp 1644511149
transform 1 0 8556 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_93
timestamp 1644511149
transform 1 0 9660 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_105
timestamp 1644511149
transform 1 0 10764 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_111
timestamp 1644511149
transform 1 0 11316 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_113
timestamp 1644511149
transform 1 0 11500 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_125
timestamp 1644511149
transform 1 0 12604 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_137
timestamp 1644511149
transform 1 0 13708 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_149
timestamp 1644511149
transform 1 0 14812 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_161
timestamp 1644511149
transform 1 0 15916 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_167
timestamp 1644511149
transform 1 0 16468 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_169
timestamp 1644511149
transform 1 0 16652 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_181
timestamp 1644511149
transform 1 0 17756 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_193
timestamp 1644511149
transform 1 0 18860 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_205
timestamp 1644511149
transform 1 0 19964 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_217
timestamp 1644511149
transform 1 0 21068 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_223
timestamp 1644511149
transform 1 0 21620 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_225
timestamp 1644511149
transform 1 0 21804 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_237
timestamp 1644511149
transform 1 0 22908 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_249
timestamp 1644511149
transform 1 0 24012 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_261
timestamp 1644511149
transform 1 0 25116 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_273
timestamp 1644511149
transform 1 0 26220 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_279
timestamp 1644511149
transform 1 0 26772 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_281
timestamp 1644511149
transform 1 0 26956 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_293
timestamp 1644511149
transform 1 0 28060 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_305
timestamp 1644511149
transform 1 0 29164 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_317
timestamp 1644511149
transform 1 0 30268 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_329
timestamp 1644511149
transform 1 0 31372 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_335
timestamp 1644511149
transform 1 0 31924 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_337
timestamp 1644511149
transform 1 0 32108 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_349
timestamp 1644511149
transform 1 0 33212 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_361
timestamp 1644511149
transform 1 0 34316 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_373
timestamp 1644511149
transform 1 0 35420 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_385
timestamp 1644511149
transform 1 0 36524 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_391
timestamp 1644511149
transform 1 0 37076 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_393
timestamp 1644511149
transform 1 0 37260 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_405
timestamp 1644511149
transform 1 0 38364 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_417
timestamp 1644511149
transform 1 0 39468 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_429
timestamp 1644511149
transform 1 0 40572 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_441
timestamp 1644511149
transform 1 0 41676 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_447
timestamp 1644511149
transform 1 0 42228 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_449
timestamp 1644511149
transform 1 0 42412 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_461
timestamp 1644511149
transform 1 0 43516 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_473
timestamp 1644511149
transform 1 0 44620 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_485
timestamp 1644511149
transform 1 0 45724 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_497
timestamp 1644511149
transform 1 0 46828 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_503
timestamp 1644511149
transform 1 0 47380 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_505
timestamp 1644511149
transform 1 0 47564 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_517
timestamp 1644511149
transform 1 0 48668 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_529
timestamp 1644511149
transform 1 0 49772 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_541
timestamp 1644511149
transform 1 0 50876 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_553
timestamp 1644511149
transform 1 0 51980 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_559
timestamp 1644511149
transform 1 0 52532 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_561
timestamp 1644511149
transform 1 0 52716 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_573
timestamp 1644511149
transform 1 0 53820 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_585
timestamp 1644511149
transform 1 0 54924 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_597
timestamp 1644511149
transform 1 0 56028 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_609
timestamp 1644511149
transform 1 0 57132 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_615
timestamp 1644511149
transform 1 0 57684 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_617
timestamp 1644511149
transform 1 0 57868 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_629
timestamp 1644511149
transform 1 0 58972 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_641
timestamp 1644511149
transform 1 0 60076 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_653
timestamp 1644511149
transform 1 0 61180 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_665
timestamp 1644511149
transform 1 0 62284 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_671
timestamp 1644511149
transform 1 0 62836 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_673
timestamp 1644511149
transform 1 0 63020 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_685
timestamp 1644511149
transform 1 0 64124 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_697
timestamp 1644511149
transform 1 0 65228 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_709
timestamp 1644511149
transform 1 0 66332 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_721
timestamp 1644511149
transform 1 0 67436 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_727
timestamp 1644511149
transform 1 0 67988 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_729
timestamp 1644511149
transform 1 0 68172 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_741
timestamp 1644511149
transform 1 0 69276 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_753
timestamp 1644511149
transform 1 0 70380 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_765
timestamp 1644511149
transform 1 0 71484 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_777
timestamp 1644511149
transform 1 0 72588 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_783
timestamp 1644511149
transform 1 0 73140 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_785
timestamp 1644511149
transform 1 0 73324 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_797
timestamp 1644511149
transform 1 0 74428 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_809
timestamp 1644511149
transform 1 0 75532 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_821
timestamp 1644511149
transform 1 0 76636 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_833
timestamp 1644511149
transform 1 0 77740 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_839
timestamp 1644511149
transform 1 0 78292 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_61_841
timestamp 1644511149
transform 1 0 78476 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_3
timestamp 1644511149
transform 1 0 1380 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_15
timestamp 1644511149
transform 1 0 2484 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_27
timestamp 1644511149
transform 1 0 3588 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_29
timestamp 1644511149
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_41
timestamp 1644511149
transform 1 0 4876 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_53
timestamp 1644511149
transform 1 0 5980 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_65
timestamp 1644511149
transform 1 0 7084 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_77
timestamp 1644511149
transform 1 0 8188 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_83
timestamp 1644511149
transform 1 0 8740 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_85
timestamp 1644511149
transform 1 0 8924 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_97
timestamp 1644511149
transform 1 0 10028 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_109
timestamp 1644511149
transform 1 0 11132 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_121
timestamp 1644511149
transform 1 0 12236 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_133
timestamp 1644511149
transform 1 0 13340 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_139
timestamp 1644511149
transform 1 0 13892 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_141
timestamp 1644511149
transform 1 0 14076 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_153
timestamp 1644511149
transform 1 0 15180 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_165
timestamp 1644511149
transform 1 0 16284 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_177
timestamp 1644511149
transform 1 0 17388 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_189
timestamp 1644511149
transform 1 0 18492 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_195
timestamp 1644511149
transform 1 0 19044 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_197
timestamp 1644511149
transform 1 0 19228 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_209
timestamp 1644511149
transform 1 0 20332 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_221
timestamp 1644511149
transform 1 0 21436 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_233
timestamp 1644511149
transform 1 0 22540 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_245
timestamp 1644511149
transform 1 0 23644 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_251
timestamp 1644511149
transform 1 0 24196 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_253
timestamp 1644511149
transform 1 0 24380 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_265
timestamp 1644511149
transform 1 0 25484 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_277
timestamp 1644511149
transform 1 0 26588 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_289
timestamp 1644511149
transform 1 0 27692 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_301
timestamp 1644511149
transform 1 0 28796 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_307
timestamp 1644511149
transform 1 0 29348 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_309
timestamp 1644511149
transform 1 0 29532 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_321
timestamp 1644511149
transform 1 0 30636 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_333
timestamp 1644511149
transform 1 0 31740 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_345
timestamp 1644511149
transform 1 0 32844 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_357
timestamp 1644511149
transform 1 0 33948 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_363
timestamp 1644511149
transform 1 0 34500 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_365
timestamp 1644511149
transform 1 0 34684 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_377
timestamp 1644511149
transform 1 0 35788 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_389
timestamp 1644511149
transform 1 0 36892 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_401
timestamp 1644511149
transform 1 0 37996 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_413
timestamp 1644511149
transform 1 0 39100 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_419
timestamp 1644511149
transform 1 0 39652 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_421
timestamp 1644511149
transform 1 0 39836 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_433
timestamp 1644511149
transform 1 0 40940 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_445
timestamp 1644511149
transform 1 0 42044 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_457
timestamp 1644511149
transform 1 0 43148 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_469
timestamp 1644511149
transform 1 0 44252 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_475
timestamp 1644511149
transform 1 0 44804 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_477
timestamp 1644511149
transform 1 0 44988 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_489
timestamp 1644511149
transform 1 0 46092 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_501
timestamp 1644511149
transform 1 0 47196 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_513
timestamp 1644511149
transform 1 0 48300 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_525
timestamp 1644511149
transform 1 0 49404 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_531
timestamp 1644511149
transform 1 0 49956 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_533
timestamp 1644511149
transform 1 0 50140 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_545
timestamp 1644511149
transform 1 0 51244 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_557
timestamp 1644511149
transform 1 0 52348 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_569
timestamp 1644511149
transform 1 0 53452 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_581
timestamp 1644511149
transform 1 0 54556 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_587
timestamp 1644511149
transform 1 0 55108 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_589
timestamp 1644511149
transform 1 0 55292 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_601
timestamp 1644511149
transform 1 0 56396 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_613
timestamp 1644511149
transform 1 0 57500 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_625
timestamp 1644511149
transform 1 0 58604 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_637
timestamp 1644511149
transform 1 0 59708 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_643
timestamp 1644511149
transform 1 0 60260 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_645
timestamp 1644511149
transform 1 0 60444 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_657
timestamp 1644511149
transform 1 0 61548 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_669
timestamp 1644511149
transform 1 0 62652 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_681
timestamp 1644511149
transform 1 0 63756 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_693
timestamp 1644511149
transform 1 0 64860 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_699
timestamp 1644511149
transform 1 0 65412 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_701
timestamp 1644511149
transform 1 0 65596 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_713
timestamp 1644511149
transform 1 0 66700 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_725
timestamp 1644511149
transform 1 0 67804 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_737
timestamp 1644511149
transform 1 0 68908 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_749
timestamp 1644511149
transform 1 0 70012 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_755
timestamp 1644511149
transform 1 0 70564 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_757
timestamp 1644511149
transform 1 0 70748 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_769
timestamp 1644511149
transform 1 0 71852 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_781
timestamp 1644511149
transform 1 0 72956 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_793
timestamp 1644511149
transform 1 0 74060 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_805
timestamp 1644511149
transform 1 0 75164 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_811
timestamp 1644511149
transform 1 0 75716 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_813
timestamp 1644511149
transform 1 0 75900 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_825
timestamp 1644511149
transform 1 0 77004 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_62_833
timestamp 1644511149
transform 1 0 77740 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_838
timestamp 1644511149
transform 1 0 78200 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_63_3
timestamp 1644511149
transform 1 0 1380 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_15
timestamp 1644511149
transform 1 0 2484 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_27
timestamp 1644511149
transform 1 0 3588 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_39
timestamp 1644511149
transform 1 0 4692 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_51
timestamp 1644511149
transform 1 0 5796 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_55
timestamp 1644511149
transform 1 0 6164 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_57
timestamp 1644511149
transform 1 0 6348 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_69
timestamp 1644511149
transform 1 0 7452 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_81
timestamp 1644511149
transform 1 0 8556 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_93
timestamp 1644511149
transform 1 0 9660 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_105
timestamp 1644511149
transform 1 0 10764 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_111
timestamp 1644511149
transform 1 0 11316 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_113
timestamp 1644511149
transform 1 0 11500 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_125
timestamp 1644511149
transform 1 0 12604 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_137
timestamp 1644511149
transform 1 0 13708 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_149
timestamp 1644511149
transform 1 0 14812 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_161
timestamp 1644511149
transform 1 0 15916 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_167
timestamp 1644511149
transform 1 0 16468 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_169
timestamp 1644511149
transform 1 0 16652 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_181
timestamp 1644511149
transform 1 0 17756 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_193
timestamp 1644511149
transform 1 0 18860 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_205
timestamp 1644511149
transform 1 0 19964 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_217
timestamp 1644511149
transform 1 0 21068 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_223
timestamp 1644511149
transform 1 0 21620 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_225
timestamp 1644511149
transform 1 0 21804 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_237
timestamp 1644511149
transform 1 0 22908 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_249
timestamp 1644511149
transform 1 0 24012 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_261
timestamp 1644511149
transform 1 0 25116 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_273
timestamp 1644511149
transform 1 0 26220 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_279
timestamp 1644511149
transform 1 0 26772 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_281
timestamp 1644511149
transform 1 0 26956 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_293
timestamp 1644511149
transform 1 0 28060 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_305
timestamp 1644511149
transform 1 0 29164 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_317
timestamp 1644511149
transform 1 0 30268 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_329
timestamp 1644511149
transform 1 0 31372 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_335
timestamp 1644511149
transform 1 0 31924 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_337
timestamp 1644511149
transform 1 0 32108 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_349
timestamp 1644511149
transform 1 0 33212 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_361
timestamp 1644511149
transform 1 0 34316 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_373
timestamp 1644511149
transform 1 0 35420 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_385
timestamp 1644511149
transform 1 0 36524 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_391
timestamp 1644511149
transform 1 0 37076 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_393
timestamp 1644511149
transform 1 0 37260 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_405
timestamp 1644511149
transform 1 0 38364 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_417
timestamp 1644511149
transform 1 0 39468 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_429
timestamp 1644511149
transform 1 0 40572 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_441
timestamp 1644511149
transform 1 0 41676 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_447
timestamp 1644511149
transform 1 0 42228 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_449
timestamp 1644511149
transform 1 0 42412 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_461
timestamp 1644511149
transform 1 0 43516 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_473
timestamp 1644511149
transform 1 0 44620 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_485
timestamp 1644511149
transform 1 0 45724 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_497
timestamp 1644511149
transform 1 0 46828 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_503
timestamp 1644511149
transform 1 0 47380 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_505
timestamp 1644511149
transform 1 0 47564 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_517
timestamp 1644511149
transform 1 0 48668 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_529
timestamp 1644511149
transform 1 0 49772 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_541
timestamp 1644511149
transform 1 0 50876 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_553
timestamp 1644511149
transform 1 0 51980 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_559
timestamp 1644511149
transform 1 0 52532 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_561
timestamp 1644511149
transform 1 0 52716 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_573
timestamp 1644511149
transform 1 0 53820 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_585
timestamp 1644511149
transform 1 0 54924 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_597
timestamp 1644511149
transform 1 0 56028 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_609
timestamp 1644511149
transform 1 0 57132 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_615
timestamp 1644511149
transform 1 0 57684 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_617
timestamp 1644511149
transform 1 0 57868 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_629
timestamp 1644511149
transform 1 0 58972 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_641
timestamp 1644511149
transform 1 0 60076 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_653
timestamp 1644511149
transform 1 0 61180 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_665
timestamp 1644511149
transform 1 0 62284 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_671
timestamp 1644511149
transform 1 0 62836 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_673
timestamp 1644511149
transform 1 0 63020 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_685
timestamp 1644511149
transform 1 0 64124 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_697
timestamp 1644511149
transform 1 0 65228 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_709
timestamp 1644511149
transform 1 0 66332 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_721
timestamp 1644511149
transform 1 0 67436 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_727
timestamp 1644511149
transform 1 0 67988 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_729
timestamp 1644511149
transform 1 0 68172 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_741
timestamp 1644511149
transform 1 0 69276 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_753
timestamp 1644511149
transform 1 0 70380 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_765
timestamp 1644511149
transform 1 0 71484 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_777
timestamp 1644511149
transform 1 0 72588 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_783
timestamp 1644511149
transform 1 0 73140 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_785
timestamp 1644511149
transform 1 0 73324 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_797
timestamp 1644511149
transform 1 0 74428 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_809
timestamp 1644511149
transform 1 0 75532 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_821
timestamp 1644511149
transform 1 0 76636 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_833
timestamp 1644511149
transform 1 0 77740 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_839
timestamp 1644511149
transform 1 0 78292 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_63_841
timestamp 1644511149
transform 1 0 78476 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_3
timestamp 1644511149
transform 1 0 1380 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_15
timestamp 1644511149
transform 1 0 2484 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_27
timestamp 1644511149
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_29
timestamp 1644511149
transform 1 0 3772 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_41
timestamp 1644511149
transform 1 0 4876 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_53
timestamp 1644511149
transform 1 0 5980 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_65
timestamp 1644511149
transform 1 0 7084 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_77
timestamp 1644511149
transform 1 0 8188 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_83
timestamp 1644511149
transform 1 0 8740 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_85
timestamp 1644511149
transform 1 0 8924 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_97
timestamp 1644511149
transform 1 0 10028 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_109
timestamp 1644511149
transform 1 0 11132 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_121
timestamp 1644511149
transform 1 0 12236 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_133
timestamp 1644511149
transform 1 0 13340 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_139
timestamp 1644511149
transform 1 0 13892 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_141
timestamp 1644511149
transform 1 0 14076 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_153
timestamp 1644511149
transform 1 0 15180 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_165
timestamp 1644511149
transform 1 0 16284 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_177
timestamp 1644511149
transform 1 0 17388 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_189
timestamp 1644511149
transform 1 0 18492 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_195
timestamp 1644511149
transform 1 0 19044 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_197
timestamp 1644511149
transform 1 0 19228 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_209
timestamp 1644511149
transform 1 0 20332 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_221
timestamp 1644511149
transform 1 0 21436 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_233
timestamp 1644511149
transform 1 0 22540 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_245
timestamp 1644511149
transform 1 0 23644 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_251
timestamp 1644511149
transform 1 0 24196 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_253
timestamp 1644511149
transform 1 0 24380 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_265
timestamp 1644511149
transform 1 0 25484 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_277
timestamp 1644511149
transform 1 0 26588 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_289
timestamp 1644511149
transform 1 0 27692 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_301
timestamp 1644511149
transform 1 0 28796 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_307
timestamp 1644511149
transform 1 0 29348 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_309
timestamp 1644511149
transform 1 0 29532 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_321
timestamp 1644511149
transform 1 0 30636 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_333
timestamp 1644511149
transform 1 0 31740 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_345
timestamp 1644511149
transform 1 0 32844 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_357
timestamp 1644511149
transform 1 0 33948 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_363
timestamp 1644511149
transform 1 0 34500 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_365
timestamp 1644511149
transform 1 0 34684 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_377
timestamp 1644511149
transform 1 0 35788 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_389
timestamp 1644511149
transform 1 0 36892 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_401
timestamp 1644511149
transform 1 0 37996 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_413
timestamp 1644511149
transform 1 0 39100 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_419
timestamp 1644511149
transform 1 0 39652 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_421
timestamp 1644511149
transform 1 0 39836 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_433
timestamp 1644511149
transform 1 0 40940 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_445
timestamp 1644511149
transform 1 0 42044 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_457
timestamp 1644511149
transform 1 0 43148 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_469
timestamp 1644511149
transform 1 0 44252 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_475
timestamp 1644511149
transform 1 0 44804 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_477
timestamp 1644511149
transform 1 0 44988 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_489
timestamp 1644511149
transform 1 0 46092 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_501
timestamp 1644511149
transform 1 0 47196 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_513
timestamp 1644511149
transform 1 0 48300 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_525
timestamp 1644511149
transform 1 0 49404 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_531
timestamp 1644511149
transform 1 0 49956 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_533
timestamp 1644511149
transform 1 0 50140 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_545
timestamp 1644511149
transform 1 0 51244 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_557
timestamp 1644511149
transform 1 0 52348 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_569
timestamp 1644511149
transform 1 0 53452 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_581
timestamp 1644511149
transform 1 0 54556 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_587
timestamp 1644511149
transform 1 0 55108 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_589
timestamp 1644511149
transform 1 0 55292 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_601
timestamp 1644511149
transform 1 0 56396 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_613
timestamp 1644511149
transform 1 0 57500 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_625
timestamp 1644511149
transform 1 0 58604 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_637
timestamp 1644511149
transform 1 0 59708 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_643
timestamp 1644511149
transform 1 0 60260 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_645
timestamp 1644511149
transform 1 0 60444 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_657
timestamp 1644511149
transform 1 0 61548 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_669
timestamp 1644511149
transform 1 0 62652 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_681
timestamp 1644511149
transform 1 0 63756 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_693
timestamp 1644511149
transform 1 0 64860 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_699
timestamp 1644511149
transform 1 0 65412 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_701
timestamp 1644511149
transform 1 0 65596 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_713
timestamp 1644511149
transform 1 0 66700 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_725
timestamp 1644511149
transform 1 0 67804 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_737
timestamp 1644511149
transform 1 0 68908 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_749
timestamp 1644511149
transform 1 0 70012 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_755
timestamp 1644511149
transform 1 0 70564 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_757
timestamp 1644511149
transform 1 0 70748 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_769
timestamp 1644511149
transform 1 0 71852 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_781
timestamp 1644511149
transform 1 0 72956 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_793
timestamp 1644511149
transform 1 0 74060 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_805
timestamp 1644511149
transform 1 0 75164 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_811
timestamp 1644511149
transform 1 0 75716 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_813
timestamp 1644511149
transform 1 0 75900 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_825
timestamp 1644511149
transform 1 0 77004 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_837
timestamp 1644511149
transform 1 0 78108 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_841
timestamp 1644511149
transform 1 0 78476 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_3
timestamp 1644511149
transform 1 0 1380 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_15
timestamp 1644511149
transform 1 0 2484 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_27
timestamp 1644511149
transform 1 0 3588 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_39
timestamp 1644511149
transform 1 0 4692 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_51
timestamp 1644511149
transform 1 0 5796 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_55
timestamp 1644511149
transform 1 0 6164 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_57
timestamp 1644511149
transform 1 0 6348 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_69
timestamp 1644511149
transform 1 0 7452 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_81
timestamp 1644511149
transform 1 0 8556 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_93
timestamp 1644511149
transform 1 0 9660 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_105
timestamp 1644511149
transform 1 0 10764 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_111
timestamp 1644511149
transform 1 0 11316 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_113
timestamp 1644511149
transform 1 0 11500 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_125
timestamp 1644511149
transform 1 0 12604 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_137
timestamp 1644511149
transform 1 0 13708 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_149
timestamp 1644511149
transform 1 0 14812 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_161
timestamp 1644511149
transform 1 0 15916 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_167
timestamp 1644511149
transform 1 0 16468 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_169
timestamp 1644511149
transform 1 0 16652 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_181
timestamp 1644511149
transform 1 0 17756 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_193
timestamp 1644511149
transform 1 0 18860 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_205
timestamp 1644511149
transform 1 0 19964 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_217
timestamp 1644511149
transform 1 0 21068 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_223
timestamp 1644511149
transform 1 0 21620 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_225
timestamp 1644511149
transform 1 0 21804 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_237
timestamp 1644511149
transform 1 0 22908 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_249
timestamp 1644511149
transform 1 0 24012 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_261
timestamp 1644511149
transform 1 0 25116 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_273
timestamp 1644511149
transform 1 0 26220 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_279
timestamp 1644511149
transform 1 0 26772 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_281
timestamp 1644511149
transform 1 0 26956 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_293
timestamp 1644511149
transform 1 0 28060 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_305
timestamp 1644511149
transform 1 0 29164 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_317
timestamp 1644511149
transform 1 0 30268 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_329
timestamp 1644511149
transform 1 0 31372 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_335
timestamp 1644511149
transform 1 0 31924 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_337
timestamp 1644511149
transform 1 0 32108 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_349
timestamp 1644511149
transform 1 0 33212 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_361
timestamp 1644511149
transform 1 0 34316 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_373
timestamp 1644511149
transform 1 0 35420 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_385
timestamp 1644511149
transform 1 0 36524 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_391
timestamp 1644511149
transform 1 0 37076 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_393
timestamp 1644511149
transform 1 0 37260 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_405
timestamp 1644511149
transform 1 0 38364 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_417
timestamp 1644511149
transform 1 0 39468 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_429
timestamp 1644511149
transform 1 0 40572 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_441
timestamp 1644511149
transform 1 0 41676 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_447
timestamp 1644511149
transform 1 0 42228 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_449
timestamp 1644511149
transform 1 0 42412 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_461
timestamp 1644511149
transform 1 0 43516 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_473
timestamp 1644511149
transform 1 0 44620 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_485
timestamp 1644511149
transform 1 0 45724 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_497
timestamp 1644511149
transform 1 0 46828 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_503
timestamp 1644511149
transform 1 0 47380 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_505
timestamp 1644511149
transform 1 0 47564 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_517
timestamp 1644511149
transform 1 0 48668 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_529
timestamp 1644511149
transform 1 0 49772 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_541
timestamp 1644511149
transform 1 0 50876 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_553
timestamp 1644511149
transform 1 0 51980 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_559
timestamp 1644511149
transform 1 0 52532 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_561
timestamp 1644511149
transform 1 0 52716 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_573
timestamp 1644511149
transform 1 0 53820 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_585
timestamp 1644511149
transform 1 0 54924 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_597
timestamp 1644511149
transform 1 0 56028 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_609
timestamp 1644511149
transform 1 0 57132 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_615
timestamp 1644511149
transform 1 0 57684 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_617
timestamp 1644511149
transform 1 0 57868 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_629
timestamp 1644511149
transform 1 0 58972 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_641
timestamp 1644511149
transform 1 0 60076 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_653
timestamp 1644511149
transform 1 0 61180 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_665
timestamp 1644511149
transform 1 0 62284 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_671
timestamp 1644511149
transform 1 0 62836 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_673
timestamp 1644511149
transform 1 0 63020 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_685
timestamp 1644511149
transform 1 0 64124 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_697
timestamp 1644511149
transform 1 0 65228 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_709
timestamp 1644511149
transform 1 0 66332 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_721
timestamp 1644511149
transform 1 0 67436 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_727
timestamp 1644511149
transform 1 0 67988 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_729
timestamp 1644511149
transform 1 0 68172 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_741
timestamp 1644511149
transform 1 0 69276 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_753
timestamp 1644511149
transform 1 0 70380 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_765
timestamp 1644511149
transform 1 0 71484 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_777
timestamp 1644511149
transform 1 0 72588 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_783
timestamp 1644511149
transform 1 0 73140 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_785
timestamp 1644511149
transform 1 0 73324 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_797
timestamp 1644511149
transform 1 0 74428 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_809
timestamp 1644511149
transform 1 0 75532 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_821
timestamp 1644511149
transform 1 0 76636 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_833
timestamp 1644511149
transform 1 0 77740 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_839
timestamp 1644511149
transform 1 0 78292 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_65_841
timestamp 1644511149
transform 1 0 78476 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_3
timestamp 1644511149
transform 1 0 1380 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_15
timestamp 1644511149
transform 1 0 2484 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_66_27
timestamp 1644511149
transform 1 0 3588 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_29
timestamp 1644511149
transform 1 0 3772 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_41
timestamp 1644511149
transform 1 0 4876 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_53
timestamp 1644511149
transform 1 0 5980 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_65
timestamp 1644511149
transform 1 0 7084 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_77
timestamp 1644511149
transform 1 0 8188 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_83
timestamp 1644511149
transform 1 0 8740 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_85
timestamp 1644511149
transform 1 0 8924 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_97
timestamp 1644511149
transform 1 0 10028 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_109
timestamp 1644511149
transform 1 0 11132 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_121
timestamp 1644511149
transform 1 0 12236 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_133
timestamp 1644511149
transform 1 0 13340 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_139
timestamp 1644511149
transform 1 0 13892 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_141
timestamp 1644511149
transform 1 0 14076 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_153
timestamp 1644511149
transform 1 0 15180 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_165
timestamp 1644511149
transform 1 0 16284 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_177
timestamp 1644511149
transform 1 0 17388 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_189
timestamp 1644511149
transform 1 0 18492 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_195
timestamp 1644511149
transform 1 0 19044 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_197
timestamp 1644511149
transform 1 0 19228 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_209
timestamp 1644511149
transform 1 0 20332 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_221
timestamp 1644511149
transform 1 0 21436 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_233
timestamp 1644511149
transform 1 0 22540 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_245
timestamp 1644511149
transform 1 0 23644 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_251
timestamp 1644511149
transform 1 0 24196 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_253
timestamp 1644511149
transform 1 0 24380 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_265
timestamp 1644511149
transform 1 0 25484 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_277
timestamp 1644511149
transform 1 0 26588 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_289
timestamp 1644511149
transform 1 0 27692 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_301
timestamp 1644511149
transform 1 0 28796 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_307
timestamp 1644511149
transform 1 0 29348 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_309
timestamp 1644511149
transform 1 0 29532 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_321
timestamp 1644511149
transform 1 0 30636 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_333
timestamp 1644511149
transform 1 0 31740 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_345
timestamp 1644511149
transform 1 0 32844 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_357
timestamp 1644511149
transform 1 0 33948 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_363
timestamp 1644511149
transform 1 0 34500 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_365
timestamp 1644511149
transform 1 0 34684 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_377
timestamp 1644511149
transform 1 0 35788 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_389
timestamp 1644511149
transform 1 0 36892 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_401
timestamp 1644511149
transform 1 0 37996 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_413
timestamp 1644511149
transform 1 0 39100 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_419
timestamp 1644511149
transform 1 0 39652 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_421
timestamp 1644511149
transform 1 0 39836 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_433
timestamp 1644511149
transform 1 0 40940 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_445
timestamp 1644511149
transform 1 0 42044 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_457
timestamp 1644511149
transform 1 0 43148 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_469
timestamp 1644511149
transform 1 0 44252 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_475
timestamp 1644511149
transform 1 0 44804 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_477
timestamp 1644511149
transform 1 0 44988 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_489
timestamp 1644511149
transform 1 0 46092 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_501
timestamp 1644511149
transform 1 0 47196 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_513
timestamp 1644511149
transform 1 0 48300 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_525
timestamp 1644511149
transform 1 0 49404 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_531
timestamp 1644511149
transform 1 0 49956 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_533
timestamp 1644511149
transform 1 0 50140 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_545
timestamp 1644511149
transform 1 0 51244 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_557
timestamp 1644511149
transform 1 0 52348 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_569
timestamp 1644511149
transform 1 0 53452 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_581
timestamp 1644511149
transform 1 0 54556 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_587
timestamp 1644511149
transform 1 0 55108 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_589
timestamp 1644511149
transform 1 0 55292 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_601
timestamp 1644511149
transform 1 0 56396 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_613
timestamp 1644511149
transform 1 0 57500 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_625
timestamp 1644511149
transform 1 0 58604 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_637
timestamp 1644511149
transform 1 0 59708 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_643
timestamp 1644511149
transform 1 0 60260 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_645
timestamp 1644511149
transform 1 0 60444 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_657
timestamp 1644511149
transform 1 0 61548 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_669
timestamp 1644511149
transform 1 0 62652 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_681
timestamp 1644511149
transform 1 0 63756 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_693
timestamp 1644511149
transform 1 0 64860 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_699
timestamp 1644511149
transform 1 0 65412 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_701
timestamp 1644511149
transform 1 0 65596 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_713
timestamp 1644511149
transform 1 0 66700 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_725
timestamp 1644511149
transform 1 0 67804 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_737
timestamp 1644511149
transform 1 0 68908 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_749
timestamp 1644511149
transform 1 0 70012 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_755
timestamp 1644511149
transform 1 0 70564 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_757
timestamp 1644511149
transform 1 0 70748 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_769
timestamp 1644511149
transform 1 0 71852 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_781
timestamp 1644511149
transform 1 0 72956 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_793
timestamp 1644511149
transform 1 0 74060 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_805
timestamp 1644511149
transform 1 0 75164 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_811
timestamp 1644511149
transform 1 0 75716 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_813
timestamp 1644511149
transform 1 0 75900 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_825
timestamp 1644511149
transform 1 0 77004 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_66_837
timestamp 1644511149
transform 1 0 78108 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_66_841
timestamp 1644511149
transform 1 0 78476 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_67_3
timestamp 1644511149
transform 1 0 1380 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_67_13
timestamp 1644511149
transform 1 0 2300 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_25
timestamp 1644511149
transform 1 0 3404 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_37
timestamp 1644511149
transform 1 0 4508 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_49
timestamp 1644511149
transform 1 0 5612 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_55
timestamp 1644511149
transform 1 0 6164 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_57
timestamp 1644511149
transform 1 0 6348 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_69
timestamp 1644511149
transform 1 0 7452 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_81
timestamp 1644511149
transform 1 0 8556 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_93
timestamp 1644511149
transform 1 0 9660 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_105
timestamp 1644511149
transform 1 0 10764 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_111
timestamp 1644511149
transform 1 0 11316 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_113
timestamp 1644511149
transform 1 0 11500 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_125
timestamp 1644511149
transform 1 0 12604 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_137
timestamp 1644511149
transform 1 0 13708 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_149
timestamp 1644511149
transform 1 0 14812 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_161
timestamp 1644511149
transform 1 0 15916 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_167
timestamp 1644511149
transform 1 0 16468 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_169
timestamp 1644511149
transform 1 0 16652 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_181
timestamp 1644511149
transform 1 0 17756 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_193
timestamp 1644511149
transform 1 0 18860 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_205
timestamp 1644511149
transform 1 0 19964 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_217
timestamp 1644511149
transform 1 0 21068 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_223
timestamp 1644511149
transform 1 0 21620 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_225
timestamp 1644511149
transform 1 0 21804 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_237
timestamp 1644511149
transform 1 0 22908 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_249
timestamp 1644511149
transform 1 0 24012 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_261
timestamp 1644511149
transform 1 0 25116 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_273
timestamp 1644511149
transform 1 0 26220 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_279
timestamp 1644511149
transform 1 0 26772 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_281
timestamp 1644511149
transform 1 0 26956 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_293
timestamp 1644511149
transform 1 0 28060 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_305
timestamp 1644511149
transform 1 0 29164 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_317
timestamp 1644511149
transform 1 0 30268 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_329
timestamp 1644511149
transform 1 0 31372 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_335
timestamp 1644511149
transform 1 0 31924 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_337
timestamp 1644511149
transform 1 0 32108 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_349
timestamp 1644511149
transform 1 0 33212 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_361
timestamp 1644511149
transform 1 0 34316 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_373
timestamp 1644511149
transform 1 0 35420 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_385
timestamp 1644511149
transform 1 0 36524 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_391
timestamp 1644511149
transform 1 0 37076 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_393
timestamp 1644511149
transform 1 0 37260 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_405
timestamp 1644511149
transform 1 0 38364 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_417
timestamp 1644511149
transform 1 0 39468 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_429
timestamp 1644511149
transform 1 0 40572 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_441
timestamp 1644511149
transform 1 0 41676 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_447
timestamp 1644511149
transform 1 0 42228 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_449
timestamp 1644511149
transform 1 0 42412 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_461
timestamp 1644511149
transform 1 0 43516 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_473
timestamp 1644511149
transform 1 0 44620 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_485
timestamp 1644511149
transform 1 0 45724 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_497
timestamp 1644511149
transform 1 0 46828 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_503
timestamp 1644511149
transform 1 0 47380 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_505
timestamp 1644511149
transform 1 0 47564 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_517
timestamp 1644511149
transform 1 0 48668 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_529
timestamp 1644511149
transform 1 0 49772 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_541
timestamp 1644511149
transform 1 0 50876 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_553
timestamp 1644511149
transform 1 0 51980 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_559
timestamp 1644511149
transform 1 0 52532 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_561
timestamp 1644511149
transform 1 0 52716 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_573
timestamp 1644511149
transform 1 0 53820 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_585
timestamp 1644511149
transform 1 0 54924 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_597
timestamp 1644511149
transform 1 0 56028 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_609
timestamp 1644511149
transform 1 0 57132 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_615
timestamp 1644511149
transform 1 0 57684 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_617
timestamp 1644511149
transform 1 0 57868 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_629
timestamp 1644511149
transform 1 0 58972 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_641
timestamp 1644511149
transform 1 0 60076 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_653
timestamp 1644511149
transform 1 0 61180 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_665
timestamp 1644511149
transform 1 0 62284 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_671
timestamp 1644511149
transform 1 0 62836 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_673
timestamp 1644511149
transform 1 0 63020 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_685
timestamp 1644511149
transform 1 0 64124 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_697
timestamp 1644511149
transform 1 0 65228 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_709
timestamp 1644511149
transform 1 0 66332 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_721
timestamp 1644511149
transform 1 0 67436 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_727
timestamp 1644511149
transform 1 0 67988 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_729
timestamp 1644511149
transform 1 0 68172 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_741
timestamp 1644511149
transform 1 0 69276 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_753
timestamp 1644511149
transform 1 0 70380 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_765
timestamp 1644511149
transform 1 0 71484 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_777
timestamp 1644511149
transform 1 0 72588 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_783
timestamp 1644511149
transform 1 0 73140 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_785
timestamp 1644511149
transform 1 0 73324 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_797
timestamp 1644511149
transform 1 0 74428 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_809
timestamp 1644511149
transform 1 0 75532 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_821
timestamp 1644511149
transform 1 0 76636 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_833
timestamp 1644511149
transform 1 0 77740 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_839
timestamp 1644511149
transform 1 0 78292 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_67_841
timestamp 1644511149
transform 1 0 78476 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_3
timestamp 1644511149
transform 1 0 1380 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_15
timestamp 1644511149
transform 1 0 2484 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_68_27
timestamp 1644511149
transform 1 0 3588 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_29
timestamp 1644511149
transform 1 0 3772 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_41
timestamp 1644511149
transform 1 0 4876 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_53
timestamp 1644511149
transform 1 0 5980 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_65
timestamp 1644511149
transform 1 0 7084 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_77
timestamp 1644511149
transform 1 0 8188 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_83
timestamp 1644511149
transform 1 0 8740 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_85
timestamp 1644511149
transform 1 0 8924 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_97
timestamp 1644511149
transform 1 0 10028 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_109
timestamp 1644511149
transform 1 0 11132 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_121
timestamp 1644511149
transform 1 0 12236 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_133
timestamp 1644511149
transform 1 0 13340 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_139
timestamp 1644511149
transform 1 0 13892 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_141
timestamp 1644511149
transform 1 0 14076 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_153
timestamp 1644511149
transform 1 0 15180 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_165
timestamp 1644511149
transform 1 0 16284 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_177
timestamp 1644511149
transform 1 0 17388 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_189
timestamp 1644511149
transform 1 0 18492 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_195
timestamp 1644511149
transform 1 0 19044 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_197
timestamp 1644511149
transform 1 0 19228 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_209
timestamp 1644511149
transform 1 0 20332 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_221
timestamp 1644511149
transform 1 0 21436 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_233
timestamp 1644511149
transform 1 0 22540 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_245
timestamp 1644511149
transform 1 0 23644 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_251
timestamp 1644511149
transform 1 0 24196 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_253
timestamp 1644511149
transform 1 0 24380 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_265
timestamp 1644511149
transform 1 0 25484 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_277
timestamp 1644511149
transform 1 0 26588 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_289
timestamp 1644511149
transform 1 0 27692 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_301
timestamp 1644511149
transform 1 0 28796 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_307
timestamp 1644511149
transform 1 0 29348 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_309
timestamp 1644511149
transform 1 0 29532 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_321
timestamp 1644511149
transform 1 0 30636 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_333
timestamp 1644511149
transform 1 0 31740 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_345
timestamp 1644511149
transform 1 0 32844 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_357
timestamp 1644511149
transform 1 0 33948 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_363
timestamp 1644511149
transform 1 0 34500 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_365
timestamp 1644511149
transform 1 0 34684 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_377
timestamp 1644511149
transform 1 0 35788 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_389
timestamp 1644511149
transform 1 0 36892 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_401
timestamp 1644511149
transform 1 0 37996 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_413
timestamp 1644511149
transform 1 0 39100 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_419
timestamp 1644511149
transform 1 0 39652 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_421
timestamp 1644511149
transform 1 0 39836 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_433
timestamp 1644511149
transform 1 0 40940 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_445
timestamp 1644511149
transform 1 0 42044 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_457
timestamp 1644511149
transform 1 0 43148 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_469
timestamp 1644511149
transform 1 0 44252 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_475
timestamp 1644511149
transform 1 0 44804 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_477
timestamp 1644511149
transform 1 0 44988 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_489
timestamp 1644511149
transform 1 0 46092 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_501
timestamp 1644511149
transform 1 0 47196 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_513
timestamp 1644511149
transform 1 0 48300 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_525
timestamp 1644511149
transform 1 0 49404 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_531
timestamp 1644511149
transform 1 0 49956 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_533
timestamp 1644511149
transform 1 0 50140 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_545
timestamp 1644511149
transform 1 0 51244 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_557
timestamp 1644511149
transform 1 0 52348 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_569
timestamp 1644511149
transform 1 0 53452 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_581
timestamp 1644511149
transform 1 0 54556 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_587
timestamp 1644511149
transform 1 0 55108 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_589
timestamp 1644511149
transform 1 0 55292 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_601
timestamp 1644511149
transform 1 0 56396 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_613
timestamp 1644511149
transform 1 0 57500 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_625
timestamp 1644511149
transform 1 0 58604 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_637
timestamp 1644511149
transform 1 0 59708 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_643
timestamp 1644511149
transform 1 0 60260 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_645
timestamp 1644511149
transform 1 0 60444 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_657
timestamp 1644511149
transform 1 0 61548 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_669
timestamp 1644511149
transform 1 0 62652 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_681
timestamp 1644511149
transform 1 0 63756 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_693
timestamp 1644511149
transform 1 0 64860 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_699
timestamp 1644511149
transform 1 0 65412 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_701
timestamp 1644511149
transform 1 0 65596 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_713
timestamp 1644511149
transform 1 0 66700 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_725
timestamp 1644511149
transform 1 0 67804 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_737
timestamp 1644511149
transform 1 0 68908 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_749
timestamp 1644511149
transform 1 0 70012 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_755
timestamp 1644511149
transform 1 0 70564 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_757
timestamp 1644511149
transform 1 0 70748 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_769
timestamp 1644511149
transform 1 0 71852 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_781
timestamp 1644511149
transform 1 0 72956 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_793
timestamp 1644511149
transform 1 0 74060 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_805
timestamp 1644511149
transform 1 0 75164 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_811
timestamp 1644511149
transform 1 0 75716 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_813
timestamp 1644511149
transform 1 0 75900 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_825
timestamp 1644511149
transform 1 0 77004 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_68_837
timestamp 1644511149
transform 1 0 78108 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_68_841
timestamp 1644511149
transform 1 0 78476 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_3
timestamp 1644511149
transform 1 0 1380 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_15
timestamp 1644511149
transform 1 0 2484 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_27
timestamp 1644511149
transform 1 0 3588 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_39
timestamp 1644511149
transform 1 0 4692 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_69_51
timestamp 1644511149
transform 1 0 5796 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_55
timestamp 1644511149
transform 1 0 6164 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_57
timestamp 1644511149
transform 1 0 6348 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_69
timestamp 1644511149
transform 1 0 7452 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_81
timestamp 1644511149
transform 1 0 8556 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_93
timestamp 1644511149
transform 1 0 9660 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_105
timestamp 1644511149
transform 1 0 10764 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_111
timestamp 1644511149
transform 1 0 11316 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_113
timestamp 1644511149
transform 1 0 11500 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_125
timestamp 1644511149
transform 1 0 12604 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_137
timestamp 1644511149
transform 1 0 13708 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_149
timestamp 1644511149
transform 1 0 14812 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_161
timestamp 1644511149
transform 1 0 15916 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_167
timestamp 1644511149
transform 1 0 16468 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_169
timestamp 1644511149
transform 1 0 16652 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_181
timestamp 1644511149
transform 1 0 17756 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_193
timestamp 1644511149
transform 1 0 18860 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_205
timestamp 1644511149
transform 1 0 19964 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_217
timestamp 1644511149
transform 1 0 21068 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_223
timestamp 1644511149
transform 1 0 21620 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_225
timestamp 1644511149
transform 1 0 21804 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_237
timestamp 1644511149
transform 1 0 22908 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_249
timestamp 1644511149
transform 1 0 24012 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_261
timestamp 1644511149
transform 1 0 25116 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_273
timestamp 1644511149
transform 1 0 26220 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_279
timestamp 1644511149
transform 1 0 26772 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_281
timestamp 1644511149
transform 1 0 26956 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_293
timestamp 1644511149
transform 1 0 28060 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_305
timestamp 1644511149
transform 1 0 29164 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_317
timestamp 1644511149
transform 1 0 30268 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_329
timestamp 1644511149
transform 1 0 31372 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_335
timestamp 1644511149
transform 1 0 31924 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_337
timestamp 1644511149
transform 1 0 32108 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_349
timestamp 1644511149
transform 1 0 33212 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_361
timestamp 1644511149
transform 1 0 34316 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_373
timestamp 1644511149
transform 1 0 35420 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_385
timestamp 1644511149
transform 1 0 36524 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_391
timestamp 1644511149
transform 1 0 37076 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_393
timestamp 1644511149
transform 1 0 37260 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_405
timestamp 1644511149
transform 1 0 38364 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_417
timestamp 1644511149
transform 1 0 39468 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_429
timestamp 1644511149
transform 1 0 40572 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_441
timestamp 1644511149
transform 1 0 41676 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_447
timestamp 1644511149
transform 1 0 42228 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_449
timestamp 1644511149
transform 1 0 42412 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_461
timestamp 1644511149
transform 1 0 43516 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_473
timestamp 1644511149
transform 1 0 44620 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_485
timestamp 1644511149
transform 1 0 45724 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_497
timestamp 1644511149
transform 1 0 46828 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_503
timestamp 1644511149
transform 1 0 47380 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_505
timestamp 1644511149
transform 1 0 47564 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_517
timestamp 1644511149
transform 1 0 48668 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_529
timestamp 1644511149
transform 1 0 49772 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_541
timestamp 1644511149
transform 1 0 50876 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_553
timestamp 1644511149
transform 1 0 51980 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_559
timestamp 1644511149
transform 1 0 52532 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_561
timestamp 1644511149
transform 1 0 52716 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_573
timestamp 1644511149
transform 1 0 53820 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_585
timestamp 1644511149
transform 1 0 54924 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_597
timestamp 1644511149
transform 1 0 56028 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_609
timestamp 1644511149
transform 1 0 57132 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_615
timestamp 1644511149
transform 1 0 57684 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_617
timestamp 1644511149
transform 1 0 57868 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_629
timestamp 1644511149
transform 1 0 58972 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_641
timestamp 1644511149
transform 1 0 60076 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_653
timestamp 1644511149
transform 1 0 61180 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_665
timestamp 1644511149
transform 1 0 62284 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_671
timestamp 1644511149
transform 1 0 62836 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_673
timestamp 1644511149
transform 1 0 63020 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_685
timestamp 1644511149
transform 1 0 64124 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_697
timestamp 1644511149
transform 1 0 65228 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_709
timestamp 1644511149
transform 1 0 66332 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_721
timestamp 1644511149
transform 1 0 67436 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_727
timestamp 1644511149
transform 1 0 67988 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_729
timestamp 1644511149
transform 1 0 68172 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_741
timestamp 1644511149
transform 1 0 69276 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_753
timestamp 1644511149
transform 1 0 70380 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_765
timestamp 1644511149
transform 1 0 71484 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_777
timestamp 1644511149
transform 1 0 72588 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_783
timestamp 1644511149
transform 1 0 73140 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_785
timestamp 1644511149
transform 1 0 73324 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_797
timestamp 1644511149
transform 1 0 74428 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_809
timestamp 1644511149
transform 1 0 75532 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_69_821
timestamp 1644511149
transform 1 0 76636 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_69_829
timestamp 1644511149
transform 1 0 77372 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_69_833
timestamp 1644511149
transform 1 0 77740 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_839
timestamp 1644511149
transform 1 0 78292 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_69_841
timestamp 1644511149
transform 1 0 78476 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_3
timestamp 1644511149
transform 1 0 1380 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_15
timestamp 1644511149
transform 1 0 2484 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_70_27
timestamp 1644511149
transform 1 0 3588 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_29
timestamp 1644511149
transform 1 0 3772 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_41
timestamp 1644511149
transform 1 0 4876 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_53
timestamp 1644511149
transform 1 0 5980 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_65
timestamp 1644511149
transform 1 0 7084 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_77
timestamp 1644511149
transform 1 0 8188 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_83
timestamp 1644511149
transform 1 0 8740 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_85
timestamp 1644511149
transform 1 0 8924 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_97
timestamp 1644511149
transform 1 0 10028 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_109
timestamp 1644511149
transform 1 0 11132 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_121
timestamp 1644511149
transform 1 0 12236 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_133
timestamp 1644511149
transform 1 0 13340 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_139
timestamp 1644511149
transform 1 0 13892 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_141
timestamp 1644511149
transform 1 0 14076 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_153
timestamp 1644511149
transform 1 0 15180 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_165
timestamp 1644511149
transform 1 0 16284 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_177
timestamp 1644511149
transform 1 0 17388 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_189
timestamp 1644511149
transform 1 0 18492 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_195
timestamp 1644511149
transform 1 0 19044 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_197
timestamp 1644511149
transform 1 0 19228 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_209
timestamp 1644511149
transform 1 0 20332 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_221
timestamp 1644511149
transform 1 0 21436 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_233
timestamp 1644511149
transform 1 0 22540 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_245
timestamp 1644511149
transform 1 0 23644 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_251
timestamp 1644511149
transform 1 0 24196 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_253
timestamp 1644511149
transform 1 0 24380 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_265
timestamp 1644511149
transform 1 0 25484 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_277
timestamp 1644511149
transform 1 0 26588 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_289
timestamp 1644511149
transform 1 0 27692 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_301
timestamp 1644511149
transform 1 0 28796 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_307
timestamp 1644511149
transform 1 0 29348 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_309
timestamp 1644511149
transform 1 0 29532 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_321
timestamp 1644511149
transform 1 0 30636 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_333
timestamp 1644511149
transform 1 0 31740 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_345
timestamp 1644511149
transform 1 0 32844 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_357
timestamp 1644511149
transform 1 0 33948 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_363
timestamp 1644511149
transform 1 0 34500 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_365
timestamp 1644511149
transform 1 0 34684 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_377
timestamp 1644511149
transform 1 0 35788 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_389
timestamp 1644511149
transform 1 0 36892 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_401
timestamp 1644511149
transform 1 0 37996 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_413
timestamp 1644511149
transform 1 0 39100 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_419
timestamp 1644511149
transform 1 0 39652 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_421
timestamp 1644511149
transform 1 0 39836 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_433
timestamp 1644511149
transform 1 0 40940 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_445
timestamp 1644511149
transform 1 0 42044 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_457
timestamp 1644511149
transform 1 0 43148 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_469
timestamp 1644511149
transform 1 0 44252 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_475
timestamp 1644511149
transform 1 0 44804 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_477
timestamp 1644511149
transform 1 0 44988 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_489
timestamp 1644511149
transform 1 0 46092 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_501
timestamp 1644511149
transform 1 0 47196 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_513
timestamp 1644511149
transform 1 0 48300 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_525
timestamp 1644511149
transform 1 0 49404 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_531
timestamp 1644511149
transform 1 0 49956 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_533
timestamp 1644511149
transform 1 0 50140 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_545
timestamp 1644511149
transform 1 0 51244 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_557
timestamp 1644511149
transform 1 0 52348 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_569
timestamp 1644511149
transform 1 0 53452 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_581
timestamp 1644511149
transform 1 0 54556 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_587
timestamp 1644511149
transform 1 0 55108 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_589
timestamp 1644511149
transform 1 0 55292 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_601
timestamp 1644511149
transform 1 0 56396 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_613
timestamp 1644511149
transform 1 0 57500 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_625
timestamp 1644511149
transform 1 0 58604 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_637
timestamp 1644511149
transform 1 0 59708 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_643
timestamp 1644511149
transform 1 0 60260 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_645
timestamp 1644511149
transform 1 0 60444 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_657
timestamp 1644511149
transform 1 0 61548 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_669
timestamp 1644511149
transform 1 0 62652 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_681
timestamp 1644511149
transform 1 0 63756 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_693
timestamp 1644511149
transform 1 0 64860 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_699
timestamp 1644511149
transform 1 0 65412 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_701
timestamp 1644511149
transform 1 0 65596 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_713
timestamp 1644511149
transform 1 0 66700 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_725
timestamp 1644511149
transform 1 0 67804 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_737
timestamp 1644511149
transform 1 0 68908 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_749
timestamp 1644511149
transform 1 0 70012 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_755
timestamp 1644511149
transform 1 0 70564 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_757
timestamp 1644511149
transform 1 0 70748 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_769
timestamp 1644511149
transform 1 0 71852 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_781
timestamp 1644511149
transform 1 0 72956 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_793
timestamp 1644511149
transform 1 0 74060 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_805
timestamp 1644511149
transform 1 0 75164 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_811
timestamp 1644511149
transform 1 0 75716 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_813
timestamp 1644511149
transform 1 0 75900 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_70_825
timestamp 1644511149
transform 1 0 77004 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_70_833
timestamp 1644511149
transform 1 0 77740 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_70_838
timestamp 1644511149
transform 1 0 78200 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_71_3
timestamp 1644511149
transform 1 0 1380 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_15
timestamp 1644511149
transform 1 0 2484 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_27
timestamp 1644511149
transform 1 0 3588 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_39
timestamp 1644511149
transform 1 0 4692 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_71_51
timestamp 1644511149
transform 1 0 5796 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_55
timestamp 1644511149
transform 1 0 6164 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_57
timestamp 1644511149
transform 1 0 6348 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_69
timestamp 1644511149
transform 1 0 7452 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_81
timestamp 1644511149
transform 1 0 8556 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_93
timestamp 1644511149
transform 1 0 9660 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_105
timestamp 1644511149
transform 1 0 10764 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_111
timestamp 1644511149
transform 1 0 11316 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_113
timestamp 1644511149
transform 1 0 11500 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_125
timestamp 1644511149
transform 1 0 12604 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_137
timestamp 1644511149
transform 1 0 13708 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_149
timestamp 1644511149
transform 1 0 14812 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_161
timestamp 1644511149
transform 1 0 15916 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_167
timestamp 1644511149
transform 1 0 16468 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_169
timestamp 1644511149
transform 1 0 16652 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_181
timestamp 1644511149
transform 1 0 17756 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_193
timestamp 1644511149
transform 1 0 18860 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_205
timestamp 1644511149
transform 1 0 19964 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_217
timestamp 1644511149
transform 1 0 21068 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_223
timestamp 1644511149
transform 1 0 21620 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_225
timestamp 1644511149
transform 1 0 21804 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_237
timestamp 1644511149
transform 1 0 22908 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_249
timestamp 1644511149
transform 1 0 24012 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_261
timestamp 1644511149
transform 1 0 25116 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_273
timestamp 1644511149
transform 1 0 26220 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_279
timestamp 1644511149
transform 1 0 26772 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_281
timestamp 1644511149
transform 1 0 26956 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_293
timestamp 1644511149
transform 1 0 28060 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_305
timestamp 1644511149
transform 1 0 29164 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_317
timestamp 1644511149
transform 1 0 30268 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_329
timestamp 1644511149
transform 1 0 31372 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_335
timestamp 1644511149
transform 1 0 31924 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_337
timestamp 1644511149
transform 1 0 32108 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_349
timestamp 1644511149
transform 1 0 33212 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_361
timestamp 1644511149
transform 1 0 34316 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_373
timestamp 1644511149
transform 1 0 35420 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_385
timestamp 1644511149
transform 1 0 36524 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_391
timestamp 1644511149
transform 1 0 37076 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_393
timestamp 1644511149
transform 1 0 37260 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_405
timestamp 1644511149
transform 1 0 38364 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_417
timestamp 1644511149
transform 1 0 39468 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_429
timestamp 1644511149
transform 1 0 40572 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_441
timestamp 1644511149
transform 1 0 41676 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_447
timestamp 1644511149
transform 1 0 42228 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_449
timestamp 1644511149
transform 1 0 42412 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_461
timestamp 1644511149
transform 1 0 43516 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_473
timestamp 1644511149
transform 1 0 44620 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_485
timestamp 1644511149
transform 1 0 45724 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_497
timestamp 1644511149
transform 1 0 46828 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_503
timestamp 1644511149
transform 1 0 47380 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_505
timestamp 1644511149
transform 1 0 47564 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_517
timestamp 1644511149
transform 1 0 48668 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_529
timestamp 1644511149
transform 1 0 49772 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_541
timestamp 1644511149
transform 1 0 50876 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_553
timestamp 1644511149
transform 1 0 51980 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_559
timestamp 1644511149
transform 1 0 52532 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_561
timestamp 1644511149
transform 1 0 52716 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_573
timestamp 1644511149
transform 1 0 53820 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_585
timestamp 1644511149
transform 1 0 54924 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_597
timestamp 1644511149
transform 1 0 56028 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_609
timestamp 1644511149
transform 1 0 57132 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_615
timestamp 1644511149
transform 1 0 57684 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_617
timestamp 1644511149
transform 1 0 57868 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_629
timestamp 1644511149
transform 1 0 58972 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_641
timestamp 1644511149
transform 1 0 60076 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_653
timestamp 1644511149
transform 1 0 61180 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_665
timestamp 1644511149
transform 1 0 62284 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_671
timestamp 1644511149
transform 1 0 62836 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_673
timestamp 1644511149
transform 1 0 63020 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_685
timestamp 1644511149
transform 1 0 64124 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_697
timestamp 1644511149
transform 1 0 65228 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_709
timestamp 1644511149
transform 1 0 66332 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_721
timestamp 1644511149
transform 1 0 67436 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_727
timestamp 1644511149
transform 1 0 67988 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_729
timestamp 1644511149
transform 1 0 68172 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_741
timestamp 1644511149
transform 1 0 69276 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_753
timestamp 1644511149
transform 1 0 70380 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_765
timestamp 1644511149
transform 1 0 71484 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_777
timestamp 1644511149
transform 1 0 72588 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_783
timestamp 1644511149
transform 1 0 73140 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_785
timestamp 1644511149
transform 1 0 73324 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_797
timestamp 1644511149
transform 1 0 74428 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_809
timestamp 1644511149
transform 1 0 75532 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_821
timestamp 1644511149
transform 1 0 76636 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_833
timestamp 1644511149
transform 1 0 77740 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_839
timestamp 1644511149
transform 1 0 78292 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_71_841
timestamp 1644511149
transform 1 0 78476 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_3
timestamp 1644511149
transform 1 0 1380 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_15
timestamp 1644511149
transform 1 0 2484 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_72_27
timestamp 1644511149
transform 1 0 3588 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_29
timestamp 1644511149
transform 1 0 3772 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_41
timestamp 1644511149
transform 1 0 4876 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_53
timestamp 1644511149
transform 1 0 5980 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_65
timestamp 1644511149
transform 1 0 7084 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_77
timestamp 1644511149
transform 1 0 8188 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_83
timestamp 1644511149
transform 1 0 8740 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_85
timestamp 1644511149
transform 1 0 8924 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_97
timestamp 1644511149
transform 1 0 10028 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_109
timestamp 1644511149
transform 1 0 11132 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_121
timestamp 1644511149
transform 1 0 12236 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_133
timestamp 1644511149
transform 1 0 13340 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_139
timestamp 1644511149
transform 1 0 13892 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_141
timestamp 1644511149
transform 1 0 14076 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_153
timestamp 1644511149
transform 1 0 15180 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_165
timestamp 1644511149
transform 1 0 16284 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_177
timestamp 1644511149
transform 1 0 17388 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_189
timestamp 1644511149
transform 1 0 18492 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_195
timestamp 1644511149
transform 1 0 19044 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_197
timestamp 1644511149
transform 1 0 19228 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_209
timestamp 1644511149
transform 1 0 20332 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_221
timestamp 1644511149
transform 1 0 21436 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_233
timestamp 1644511149
transform 1 0 22540 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_245
timestamp 1644511149
transform 1 0 23644 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_251
timestamp 1644511149
transform 1 0 24196 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_253
timestamp 1644511149
transform 1 0 24380 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_265
timestamp 1644511149
transform 1 0 25484 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_277
timestamp 1644511149
transform 1 0 26588 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_289
timestamp 1644511149
transform 1 0 27692 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_301
timestamp 1644511149
transform 1 0 28796 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_307
timestamp 1644511149
transform 1 0 29348 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_309
timestamp 1644511149
transform 1 0 29532 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_321
timestamp 1644511149
transform 1 0 30636 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_333
timestamp 1644511149
transform 1 0 31740 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_345
timestamp 1644511149
transform 1 0 32844 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_357
timestamp 1644511149
transform 1 0 33948 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_363
timestamp 1644511149
transform 1 0 34500 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_365
timestamp 1644511149
transform 1 0 34684 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_377
timestamp 1644511149
transform 1 0 35788 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_389
timestamp 1644511149
transform 1 0 36892 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_401
timestamp 1644511149
transform 1 0 37996 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_413
timestamp 1644511149
transform 1 0 39100 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_419
timestamp 1644511149
transform 1 0 39652 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_421
timestamp 1644511149
transform 1 0 39836 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_433
timestamp 1644511149
transform 1 0 40940 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_445
timestamp 1644511149
transform 1 0 42044 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_457
timestamp 1644511149
transform 1 0 43148 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_469
timestamp 1644511149
transform 1 0 44252 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_475
timestamp 1644511149
transform 1 0 44804 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_477
timestamp 1644511149
transform 1 0 44988 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_489
timestamp 1644511149
transform 1 0 46092 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_501
timestamp 1644511149
transform 1 0 47196 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_513
timestamp 1644511149
transform 1 0 48300 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_525
timestamp 1644511149
transform 1 0 49404 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_531
timestamp 1644511149
transform 1 0 49956 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_533
timestamp 1644511149
transform 1 0 50140 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_545
timestamp 1644511149
transform 1 0 51244 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_557
timestamp 1644511149
transform 1 0 52348 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_569
timestamp 1644511149
transform 1 0 53452 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_581
timestamp 1644511149
transform 1 0 54556 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_587
timestamp 1644511149
transform 1 0 55108 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_589
timestamp 1644511149
transform 1 0 55292 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_601
timestamp 1644511149
transform 1 0 56396 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_613
timestamp 1644511149
transform 1 0 57500 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_625
timestamp 1644511149
transform 1 0 58604 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_637
timestamp 1644511149
transform 1 0 59708 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_643
timestamp 1644511149
transform 1 0 60260 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_645
timestamp 1644511149
transform 1 0 60444 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_657
timestamp 1644511149
transform 1 0 61548 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_669
timestamp 1644511149
transform 1 0 62652 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_681
timestamp 1644511149
transform 1 0 63756 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_693
timestamp 1644511149
transform 1 0 64860 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_699
timestamp 1644511149
transform 1 0 65412 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_701
timestamp 1644511149
transform 1 0 65596 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_713
timestamp 1644511149
transform 1 0 66700 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_725
timestamp 1644511149
transform 1 0 67804 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_737
timestamp 1644511149
transform 1 0 68908 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_749
timestamp 1644511149
transform 1 0 70012 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_755
timestamp 1644511149
transform 1 0 70564 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_757
timestamp 1644511149
transform 1 0 70748 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_769
timestamp 1644511149
transform 1 0 71852 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_781
timestamp 1644511149
transform 1 0 72956 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_793
timestamp 1644511149
transform 1 0 74060 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_805
timestamp 1644511149
transform 1 0 75164 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_811
timestamp 1644511149
transform 1 0 75716 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_813
timestamp 1644511149
transform 1 0 75900 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_825
timestamp 1644511149
transform 1 0 77004 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_72_837
timestamp 1644511149
transform 1 0 78108 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_72_841
timestamp 1644511149
transform 1 0 78476 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_3
timestamp 1644511149
transform 1 0 1380 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_15
timestamp 1644511149
transform 1 0 2484 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_27
timestamp 1644511149
transform 1 0 3588 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_39
timestamp 1644511149
transform 1 0 4692 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_73_51
timestamp 1644511149
transform 1 0 5796 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_55
timestamp 1644511149
transform 1 0 6164 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_57
timestamp 1644511149
transform 1 0 6348 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_69
timestamp 1644511149
transform 1 0 7452 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_81
timestamp 1644511149
transform 1 0 8556 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_93
timestamp 1644511149
transform 1 0 9660 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_105
timestamp 1644511149
transform 1 0 10764 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_111
timestamp 1644511149
transform 1 0 11316 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_113
timestamp 1644511149
transform 1 0 11500 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_125
timestamp 1644511149
transform 1 0 12604 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_137
timestamp 1644511149
transform 1 0 13708 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_149
timestamp 1644511149
transform 1 0 14812 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_161
timestamp 1644511149
transform 1 0 15916 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_167
timestamp 1644511149
transform 1 0 16468 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_169
timestamp 1644511149
transform 1 0 16652 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_181
timestamp 1644511149
transform 1 0 17756 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_193
timestamp 1644511149
transform 1 0 18860 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_205
timestamp 1644511149
transform 1 0 19964 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_217
timestamp 1644511149
transform 1 0 21068 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_223
timestamp 1644511149
transform 1 0 21620 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_225
timestamp 1644511149
transform 1 0 21804 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_237
timestamp 1644511149
transform 1 0 22908 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_249
timestamp 1644511149
transform 1 0 24012 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_261
timestamp 1644511149
transform 1 0 25116 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_273
timestamp 1644511149
transform 1 0 26220 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_279
timestamp 1644511149
transform 1 0 26772 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_281
timestamp 1644511149
transform 1 0 26956 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_293
timestamp 1644511149
transform 1 0 28060 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_305
timestamp 1644511149
transform 1 0 29164 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_317
timestamp 1644511149
transform 1 0 30268 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_329
timestamp 1644511149
transform 1 0 31372 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_335
timestamp 1644511149
transform 1 0 31924 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_337
timestamp 1644511149
transform 1 0 32108 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_349
timestamp 1644511149
transform 1 0 33212 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_361
timestamp 1644511149
transform 1 0 34316 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_373
timestamp 1644511149
transform 1 0 35420 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_385
timestamp 1644511149
transform 1 0 36524 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_391
timestamp 1644511149
transform 1 0 37076 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_393
timestamp 1644511149
transform 1 0 37260 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_405
timestamp 1644511149
transform 1 0 38364 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_417
timestamp 1644511149
transform 1 0 39468 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_429
timestamp 1644511149
transform 1 0 40572 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_441
timestamp 1644511149
transform 1 0 41676 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_447
timestamp 1644511149
transform 1 0 42228 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_449
timestamp 1644511149
transform 1 0 42412 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_461
timestamp 1644511149
transform 1 0 43516 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_473
timestamp 1644511149
transform 1 0 44620 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_485
timestamp 1644511149
transform 1 0 45724 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_497
timestamp 1644511149
transform 1 0 46828 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_503
timestamp 1644511149
transform 1 0 47380 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_505
timestamp 1644511149
transform 1 0 47564 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_517
timestamp 1644511149
transform 1 0 48668 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_529
timestamp 1644511149
transform 1 0 49772 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_541
timestamp 1644511149
transform 1 0 50876 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_553
timestamp 1644511149
transform 1 0 51980 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_559
timestamp 1644511149
transform 1 0 52532 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_561
timestamp 1644511149
transform 1 0 52716 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_573
timestamp 1644511149
transform 1 0 53820 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_585
timestamp 1644511149
transform 1 0 54924 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_597
timestamp 1644511149
transform 1 0 56028 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_609
timestamp 1644511149
transform 1 0 57132 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_615
timestamp 1644511149
transform 1 0 57684 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_617
timestamp 1644511149
transform 1 0 57868 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_629
timestamp 1644511149
transform 1 0 58972 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_641
timestamp 1644511149
transform 1 0 60076 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_653
timestamp 1644511149
transform 1 0 61180 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_665
timestamp 1644511149
transform 1 0 62284 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_671
timestamp 1644511149
transform 1 0 62836 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_673
timestamp 1644511149
transform 1 0 63020 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_685
timestamp 1644511149
transform 1 0 64124 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_697
timestamp 1644511149
transform 1 0 65228 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_709
timestamp 1644511149
transform 1 0 66332 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_721
timestamp 1644511149
transform 1 0 67436 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_727
timestamp 1644511149
transform 1 0 67988 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_729
timestamp 1644511149
transform 1 0 68172 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_741
timestamp 1644511149
transform 1 0 69276 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_753
timestamp 1644511149
transform 1 0 70380 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_765
timestamp 1644511149
transform 1 0 71484 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_777
timestamp 1644511149
transform 1 0 72588 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_783
timestamp 1644511149
transform 1 0 73140 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_785
timestamp 1644511149
transform 1 0 73324 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_797
timestamp 1644511149
transform 1 0 74428 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_809
timestamp 1644511149
transform 1 0 75532 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_821
timestamp 1644511149
transform 1 0 76636 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_833
timestamp 1644511149
transform 1 0 77740 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_839
timestamp 1644511149
transform 1 0 78292 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_73_841
timestamp 1644511149
transform 1 0 78476 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_3
timestamp 1644511149
transform 1 0 1380 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_15
timestamp 1644511149
transform 1 0 2484 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_74_27
timestamp 1644511149
transform 1 0 3588 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_29
timestamp 1644511149
transform 1 0 3772 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_41
timestamp 1644511149
transform 1 0 4876 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_53
timestamp 1644511149
transform 1 0 5980 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_65
timestamp 1644511149
transform 1 0 7084 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_77
timestamp 1644511149
transform 1 0 8188 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_83
timestamp 1644511149
transform 1 0 8740 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_85
timestamp 1644511149
transform 1 0 8924 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_97
timestamp 1644511149
transform 1 0 10028 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_109
timestamp 1644511149
transform 1 0 11132 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_121
timestamp 1644511149
transform 1 0 12236 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_133
timestamp 1644511149
transform 1 0 13340 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_139
timestamp 1644511149
transform 1 0 13892 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_141
timestamp 1644511149
transform 1 0 14076 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_153
timestamp 1644511149
transform 1 0 15180 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_165
timestamp 1644511149
transform 1 0 16284 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_177
timestamp 1644511149
transform 1 0 17388 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_189
timestamp 1644511149
transform 1 0 18492 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_195
timestamp 1644511149
transform 1 0 19044 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_197
timestamp 1644511149
transform 1 0 19228 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_209
timestamp 1644511149
transform 1 0 20332 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_221
timestamp 1644511149
transform 1 0 21436 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_233
timestamp 1644511149
transform 1 0 22540 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_245
timestamp 1644511149
transform 1 0 23644 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_251
timestamp 1644511149
transform 1 0 24196 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_253
timestamp 1644511149
transform 1 0 24380 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_265
timestamp 1644511149
transform 1 0 25484 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_277
timestamp 1644511149
transform 1 0 26588 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_289
timestamp 1644511149
transform 1 0 27692 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_301
timestamp 1644511149
transform 1 0 28796 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_307
timestamp 1644511149
transform 1 0 29348 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_309
timestamp 1644511149
transform 1 0 29532 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_321
timestamp 1644511149
transform 1 0 30636 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_333
timestamp 1644511149
transform 1 0 31740 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_345
timestamp 1644511149
transform 1 0 32844 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_357
timestamp 1644511149
transform 1 0 33948 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_363
timestamp 1644511149
transform 1 0 34500 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_365
timestamp 1644511149
transform 1 0 34684 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_377
timestamp 1644511149
transform 1 0 35788 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_389
timestamp 1644511149
transform 1 0 36892 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_401
timestamp 1644511149
transform 1 0 37996 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_413
timestamp 1644511149
transform 1 0 39100 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_419
timestamp 1644511149
transform 1 0 39652 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_421
timestamp 1644511149
transform 1 0 39836 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_433
timestamp 1644511149
transform 1 0 40940 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_445
timestamp 1644511149
transform 1 0 42044 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_457
timestamp 1644511149
transform 1 0 43148 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_469
timestamp 1644511149
transform 1 0 44252 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_475
timestamp 1644511149
transform 1 0 44804 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_477
timestamp 1644511149
transform 1 0 44988 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_489
timestamp 1644511149
transform 1 0 46092 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_501
timestamp 1644511149
transform 1 0 47196 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_513
timestamp 1644511149
transform 1 0 48300 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_525
timestamp 1644511149
transform 1 0 49404 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_531
timestamp 1644511149
transform 1 0 49956 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_533
timestamp 1644511149
transform 1 0 50140 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_545
timestamp 1644511149
transform 1 0 51244 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_557
timestamp 1644511149
transform 1 0 52348 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_569
timestamp 1644511149
transform 1 0 53452 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_581
timestamp 1644511149
transform 1 0 54556 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_587
timestamp 1644511149
transform 1 0 55108 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_589
timestamp 1644511149
transform 1 0 55292 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_601
timestamp 1644511149
transform 1 0 56396 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_613
timestamp 1644511149
transform 1 0 57500 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_625
timestamp 1644511149
transform 1 0 58604 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_637
timestamp 1644511149
transform 1 0 59708 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_643
timestamp 1644511149
transform 1 0 60260 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_645
timestamp 1644511149
transform 1 0 60444 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_657
timestamp 1644511149
transform 1 0 61548 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_669
timestamp 1644511149
transform 1 0 62652 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_681
timestamp 1644511149
transform 1 0 63756 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_693
timestamp 1644511149
transform 1 0 64860 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_699
timestamp 1644511149
transform 1 0 65412 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_701
timestamp 1644511149
transform 1 0 65596 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_713
timestamp 1644511149
transform 1 0 66700 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_725
timestamp 1644511149
transform 1 0 67804 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_737
timestamp 1644511149
transform 1 0 68908 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_749
timestamp 1644511149
transform 1 0 70012 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_755
timestamp 1644511149
transform 1 0 70564 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_757
timestamp 1644511149
transform 1 0 70748 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_769
timestamp 1644511149
transform 1 0 71852 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_781
timestamp 1644511149
transform 1 0 72956 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_793
timestamp 1644511149
transform 1 0 74060 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_805
timestamp 1644511149
transform 1 0 75164 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_811
timestamp 1644511149
transform 1 0 75716 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_813
timestamp 1644511149
transform 1 0 75900 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_74_825
timestamp 1644511149
transform 1 0 77004 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_74_829
timestamp 1644511149
transform 1 0 77372 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_74_834
timestamp 1644511149
transform 1 0 77832 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_75_3
timestamp 1644511149
transform 1 0 1380 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_75_13
timestamp 1644511149
transform 1 0 2300 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_25
timestamp 1644511149
transform 1 0 3404 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_37
timestamp 1644511149
transform 1 0 4508 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_49
timestamp 1644511149
transform 1 0 5612 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_55
timestamp 1644511149
transform 1 0 6164 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_57
timestamp 1644511149
transform 1 0 6348 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_69
timestamp 1644511149
transform 1 0 7452 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_81
timestamp 1644511149
transform 1 0 8556 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_93
timestamp 1644511149
transform 1 0 9660 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_105
timestamp 1644511149
transform 1 0 10764 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_111
timestamp 1644511149
transform 1 0 11316 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_113
timestamp 1644511149
transform 1 0 11500 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_125
timestamp 1644511149
transform 1 0 12604 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_137
timestamp 1644511149
transform 1 0 13708 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_149
timestamp 1644511149
transform 1 0 14812 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_161
timestamp 1644511149
transform 1 0 15916 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_167
timestamp 1644511149
transform 1 0 16468 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_169
timestamp 1644511149
transform 1 0 16652 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_181
timestamp 1644511149
transform 1 0 17756 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_193
timestamp 1644511149
transform 1 0 18860 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_205
timestamp 1644511149
transform 1 0 19964 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_217
timestamp 1644511149
transform 1 0 21068 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_223
timestamp 1644511149
transform 1 0 21620 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_225
timestamp 1644511149
transform 1 0 21804 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_237
timestamp 1644511149
transform 1 0 22908 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_249
timestamp 1644511149
transform 1 0 24012 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_261
timestamp 1644511149
transform 1 0 25116 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_273
timestamp 1644511149
transform 1 0 26220 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_279
timestamp 1644511149
transform 1 0 26772 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_281
timestamp 1644511149
transform 1 0 26956 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_293
timestamp 1644511149
transform 1 0 28060 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_305
timestamp 1644511149
transform 1 0 29164 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_317
timestamp 1644511149
transform 1 0 30268 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_329
timestamp 1644511149
transform 1 0 31372 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_335
timestamp 1644511149
transform 1 0 31924 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_337
timestamp 1644511149
transform 1 0 32108 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_349
timestamp 1644511149
transform 1 0 33212 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_361
timestamp 1644511149
transform 1 0 34316 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_373
timestamp 1644511149
transform 1 0 35420 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_385
timestamp 1644511149
transform 1 0 36524 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_391
timestamp 1644511149
transform 1 0 37076 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_393
timestamp 1644511149
transform 1 0 37260 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_405
timestamp 1644511149
transform 1 0 38364 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_417
timestamp 1644511149
transform 1 0 39468 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_429
timestamp 1644511149
transform 1 0 40572 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_441
timestamp 1644511149
transform 1 0 41676 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_447
timestamp 1644511149
transform 1 0 42228 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_449
timestamp 1644511149
transform 1 0 42412 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_461
timestamp 1644511149
transform 1 0 43516 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_473
timestamp 1644511149
transform 1 0 44620 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_485
timestamp 1644511149
transform 1 0 45724 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_497
timestamp 1644511149
transform 1 0 46828 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_503
timestamp 1644511149
transform 1 0 47380 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_505
timestamp 1644511149
transform 1 0 47564 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_517
timestamp 1644511149
transform 1 0 48668 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_529
timestamp 1644511149
transform 1 0 49772 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_541
timestamp 1644511149
transform 1 0 50876 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_553
timestamp 1644511149
transform 1 0 51980 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_559
timestamp 1644511149
transform 1 0 52532 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_561
timestamp 1644511149
transform 1 0 52716 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_573
timestamp 1644511149
transform 1 0 53820 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_585
timestamp 1644511149
transform 1 0 54924 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_597
timestamp 1644511149
transform 1 0 56028 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_609
timestamp 1644511149
transform 1 0 57132 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_615
timestamp 1644511149
transform 1 0 57684 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_617
timestamp 1644511149
transform 1 0 57868 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_629
timestamp 1644511149
transform 1 0 58972 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_641
timestamp 1644511149
transform 1 0 60076 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_653
timestamp 1644511149
transform 1 0 61180 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_665
timestamp 1644511149
transform 1 0 62284 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_671
timestamp 1644511149
transform 1 0 62836 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_673
timestamp 1644511149
transform 1 0 63020 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_685
timestamp 1644511149
transform 1 0 64124 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_697
timestamp 1644511149
transform 1 0 65228 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_709
timestamp 1644511149
transform 1 0 66332 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_721
timestamp 1644511149
transform 1 0 67436 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_727
timestamp 1644511149
transform 1 0 67988 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_729
timestamp 1644511149
transform 1 0 68172 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_741
timestamp 1644511149
transform 1 0 69276 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_753
timestamp 1644511149
transform 1 0 70380 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_765
timestamp 1644511149
transform 1 0 71484 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_777
timestamp 1644511149
transform 1 0 72588 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_783
timestamp 1644511149
transform 1 0 73140 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_785
timestamp 1644511149
transform 1 0 73324 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_797
timestamp 1644511149
transform 1 0 74428 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_809
timestamp 1644511149
transform 1 0 75532 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_821
timestamp 1644511149
transform 1 0 76636 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_833
timestamp 1644511149
transform 1 0 77740 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_839
timestamp 1644511149
transform 1 0 78292 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_75_841
timestamp 1644511149
transform 1 0 78476 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_3
timestamp 1644511149
transform 1 0 1380 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_15
timestamp 1644511149
transform 1 0 2484 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_76_27
timestamp 1644511149
transform 1 0 3588 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_29
timestamp 1644511149
transform 1 0 3772 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_41
timestamp 1644511149
transform 1 0 4876 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_53
timestamp 1644511149
transform 1 0 5980 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_65
timestamp 1644511149
transform 1 0 7084 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_77
timestamp 1644511149
transform 1 0 8188 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_83
timestamp 1644511149
transform 1 0 8740 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_85
timestamp 1644511149
transform 1 0 8924 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_97
timestamp 1644511149
transform 1 0 10028 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_109
timestamp 1644511149
transform 1 0 11132 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_121
timestamp 1644511149
transform 1 0 12236 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_133
timestamp 1644511149
transform 1 0 13340 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_139
timestamp 1644511149
transform 1 0 13892 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_141
timestamp 1644511149
transform 1 0 14076 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_153
timestamp 1644511149
transform 1 0 15180 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_165
timestamp 1644511149
transform 1 0 16284 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_177
timestamp 1644511149
transform 1 0 17388 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_189
timestamp 1644511149
transform 1 0 18492 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_195
timestamp 1644511149
transform 1 0 19044 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_197
timestamp 1644511149
transform 1 0 19228 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_209
timestamp 1644511149
transform 1 0 20332 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_221
timestamp 1644511149
transform 1 0 21436 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_233
timestamp 1644511149
transform 1 0 22540 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_245
timestamp 1644511149
transform 1 0 23644 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_251
timestamp 1644511149
transform 1 0 24196 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_253
timestamp 1644511149
transform 1 0 24380 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_265
timestamp 1644511149
transform 1 0 25484 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_277
timestamp 1644511149
transform 1 0 26588 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_289
timestamp 1644511149
transform 1 0 27692 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_301
timestamp 1644511149
transform 1 0 28796 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_307
timestamp 1644511149
transform 1 0 29348 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_309
timestamp 1644511149
transform 1 0 29532 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_321
timestamp 1644511149
transform 1 0 30636 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_333
timestamp 1644511149
transform 1 0 31740 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_345
timestamp 1644511149
transform 1 0 32844 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_357
timestamp 1644511149
transform 1 0 33948 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_363
timestamp 1644511149
transform 1 0 34500 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_365
timestamp 1644511149
transform 1 0 34684 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_377
timestamp 1644511149
transform 1 0 35788 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_389
timestamp 1644511149
transform 1 0 36892 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_401
timestamp 1644511149
transform 1 0 37996 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_413
timestamp 1644511149
transform 1 0 39100 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_419
timestamp 1644511149
transform 1 0 39652 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_421
timestamp 1644511149
transform 1 0 39836 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_433
timestamp 1644511149
transform 1 0 40940 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_445
timestamp 1644511149
transform 1 0 42044 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_457
timestamp 1644511149
transform 1 0 43148 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_469
timestamp 1644511149
transform 1 0 44252 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_475
timestamp 1644511149
transform 1 0 44804 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_477
timestamp 1644511149
transform 1 0 44988 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_489
timestamp 1644511149
transform 1 0 46092 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_501
timestamp 1644511149
transform 1 0 47196 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_513
timestamp 1644511149
transform 1 0 48300 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_525
timestamp 1644511149
transform 1 0 49404 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_531
timestamp 1644511149
transform 1 0 49956 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_533
timestamp 1644511149
transform 1 0 50140 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_545
timestamp 1644511149
transform 1 0 51244 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_557
timestamp 1644511149
transform 1 0 52348 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_569
timestamp 1644511149
transform 1 0 53452 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_581
timestamp 1644511149
transform 1 0 54556 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_587
timestamp 1644511149
transform 1 0 55108 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_589
timestamp 1644511149
transform 1 0 55292 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_601
timestamp 1644511149
transform 1 0 56396 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_613
timestamp 1644511149
transform 1 0 57500 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_625
timestamp 1644511149
transform 1 0 58604 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_637
timestamp 1644511149
transform 1 0 59708 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_643
timestamp 1644511149
transform 1 0 60260 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_645
timestamp 1644511149
transform 1 0 60444 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_657
timestamp 1644511149
transform 1 0 61548 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_669
timestamp 1644511149
transform 1 0 62652 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_681
timestamp 1644511149
transform 1 0 63756 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_693
timestamp 1644511149
transform 1 0 64860 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_699
timestamp 1644511149
transform 1 0 65412 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_701
timestamp 1644511149
transform 1 0 65596 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_713
timestamp 1644511149
transform 1 0 66700 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_725
timestamp 1644511149
transform 1 0 67804 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_737
timestamp 1644511149
transform 1 0 68908 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_749
timestamp 1644511149
transform 1 0 70012 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_755
timestamp 1644511149
transform 1 0 70564 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_757
timestamp 1644511149
transform 1 0 70748 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_769
timestamp 1644511149
transform 1 0 71852 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_781
timestamp 1644511149
transform 1 0 72956 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_793
timestamp 1644511149
transform 1 0 74060 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_805
timestamp 1644511149
transform 1 0 75164 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_811
timestamp 1644511149
transform 1 0 75716 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_813
timestamp 1644511149
transform 1 0 75900 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_76_825
timestamp 1644511149
transform 1 0 77004 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_76_833
timestamp 1644511149
transform 1 0 77740 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_76_838
timestamp 1644511149
transform 1 0 78200 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_77_3
timestamp 1644511149
transform 1 0 1380 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_15
timestamp 1644511149
transform 1 0 2484 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_27
timestamp 1644511149
transform 1 0 3588 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_39
timestamp 1644511149
transform 1 0 4692 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_77_51
timestamp 1644511149
transform 1 0 5796 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_55
timestamp 1644511149
transform 1 0 6164 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_57
timestamp 1644511149
transform 1 0 6348 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_69
timestamp 1644511149
transform 1 0 7452 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_81
timestamp 1644511149
transform 1 0 8556 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_93
timestamp 1644511149
transform 1 0 9660 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_105
timestamp 1644511149
transform 1 0 10764 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_111
timestamp 1644511149
transform 1 0 11316 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_113
timestamp 1644511149
transform 1 0 11500 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_125
timestamp 1644511149
transform 1 0 12604 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_137
timestamp 1644511149
transform 1 0 13708 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_149
timestamp 1644511149
transform 1 0 14812 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_161
timestamp 1644511149
transform 1 0 15916 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_167
timestamp 1644511149
transform 1 0 16468 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_169
timestamp 1644511149
transform 1 0 16652 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_181
timestamp 1644511149
transform 1 0 17756 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_193
timestamp 1644511149
transform 1 0 18860 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_205
timestamp 1644511149
transform 1 0 19964 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_217
timestamp 1644511149
transform 1 0 21068 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_223
timestamp 1644511149
transform 1 0 21620 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_225
timestamp 1644511149
transform 1 0 21804 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_237
timestamp 1644511149
transform 1 0 22908 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_249
timestamp 1644511149
transform 1 0 24012 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_261
timestamp 1644511149
transform 1 0 25116 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_273
timestamp 1644511149
transform 1 0 26220 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_279
timestamp 1644511149
transform 1 0 26772 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_281
timestamp 1644511149
transform 1 0 26956 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_293
timestamp 1644511149
transform 1 0 28060 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_305
timestamp 1644511149
transform 1 0 29164 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_317
timestamp 1644511149
transform 1 0 30268 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_329
timestamp 1644511149
transform 1 0 31372 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_335
timestamp 1644511149
transform 1 0 31924 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_337
timestamp 1644511149
transform 1 0 32108 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_349
timestamp 1644511149
transform 1 0 33212 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_361
timestamp 1644511149
transform 1 0 34316 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_373
timestamp 1644511149
transform 1 0 35420 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_385
timestamp 1644511149
transform 1 0 36524 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_391
timestamp 1644511149
transform 1 0 37076 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_393
timestamp 1644511149
transform 1 0 37260 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_405
timestamp 1644511149
transform 1 0 38364 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_417
timestamp 1644511149
transform 1 0 39468 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_429
timestamp 1644511149
transform 1 0 40572 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_441
timestamp 1644511149
transform 1 0 41676 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_447
timestamp 1644511149
transform 1 0 42228 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_449
timestamp 1644511149
transform 1 0 42412 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_461
timestamp 1644511149
transform 1 0 43516 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_473
timestamp 1644511149
transform 1 0 44620 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_485
timestamp 1644511149
transform 1 0 45724 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_497
timestamp 1644511149
transform 1 0 46828 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_503
timestamp 1644511149
transform 1 0 47380 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_505
timestamp 1644511149
transform 1 0 47564 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_517
timestamp 1644511149
transform 1 0 48668 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_529
timestamp 1644511149
transform 1 0 49772 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_541
timestamp 1644511149
transform 1 0 50876 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_553
timestamp 1644511149
transform 1 0 51980 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_559
timestamp 1644511149
transform 1 0 52532 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_561
timestamp 1644511149
transform 1 0 52716 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_573
timestamp 1644511149
transform 1 0 53820 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_585
timestamp 1644511149
transform 1 0 54924 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_597
timestamp 1644511149
transform 1 0 56028 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_609
timestamp 1644511149
transform 1 0 57132 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_615
timestamp 1644511149
transform 1 0 57684 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_617
timestamp 1644511149
transform 1 0 57868 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_629
timestamp 1644511149
transform 1 0 58972 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_641
timestamp 1644511149
transform 1 0 60076 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_653
timestamp 1644511149
transform 1 0 61180 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_665
timestamp 1644511149
transform 1 0 62284 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_671
timestamp 1644511149
transform 1 0 62836 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_673
timestamp 1644511149
transform 1 0 63020 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_685
timestamp 1644511149
transform 1 0 64124 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_697
timestamp 1644511149
transform 1 0 65228 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_709
timestamp 1644511149
transform 1 0 66332 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_721
timestamp 1644511149
transform 1 0 67436 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_727
timestamp 1644511149
transform 1 0 67988 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_729
timestamp 1644511149
transform 1 0 68172 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_741
timestamp 1644511149
transform 1 0 69276 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_753
timestamp 1644511149
transform 1 0 70380 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_765
timestamp 1644511149
transform 1 0 71484 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_777
timestamp 1644511149
transform 1 0 72588 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_783
timestamp 1644511149
transform 1 0 73140 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_785
timestamp 1644511149
transform 1 0 73324 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_797
timestamp 1644511149
transform 1 0 74428 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_809
timestamp 1644511149
transform 1 0 75532 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_821
timestamp 1644511149
transform 1 0 76636 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_833
timestamp 1644511149
transform 1 0 77740 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_839
timestamp 1644511149
transform 1 0 78292 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_77_841
timestamp 1644511149
transform 1 0 78476 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_3
timestamp 1644511149
transform 1 0 1380 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_15
timestamp 1644511149
transform 1 0 2484 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_78_27
timestamp 1644511149
transform 1 0 3588 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_29
timestamp 1644511149
transform 1 0 3772 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_41
timestamp 1644511149
transform 1 0 4876 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_53
timestamp 1644511149
transform 1 0 5980 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_65
timestamp 1644511149
transform 1 0 7084 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_77
timestamp 1644511149
transform 1 0 8188 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_83
timestamp 1644511149
transform 1 0 8740 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_85
timestamp 1644511149
transform 1 0 8924 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_97
timestamp 1644511149
transform 1 0 10028 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_109
timestamp 1644511149
transform 1 0 11132 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_121
timestamp 1644511149
transform 1 0 12236 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_133
timestamp 1644511149
transform 1 0 13340 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_139
timestamp 1644511149
transform 1 0 13892 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_141
timestamp 1644511149
transform 1 0 14076 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_153
timestamp 1644511149
transform 1 0 15180 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_165
timestamp 1644511149
transform 1 0 16284 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_177
timestamp 1644511149
transform 1 0 17388 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_189
timestamp 1644511149
transform 1 0 18492 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_195
timestamp 1644511149
transform 1 0 19044 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_197
timestamp 1644511149
transform 1 0 19228 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_209
timestamp 1644511149
transform 1 0 20332 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_221
timestamp 1644511149
transform 1 0 21436 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_233
timestamp 1644511149
transform 1 0 22540 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_245
timestamp 1644511149
transform 1 0 23644 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_251
timestamp 1644511149
transform 1 0 24196 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_253
timestamp 1644511149
transform 1 0 24380 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_265
timestamp 1644511149
transform 1 0 25484 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_277
timestamp 1644511149
transform 1 0 26588 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_289
timestamp 1644511149
transform 1 0 27692 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_301
timestamp 1644511149
transform 1 0 28796 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_307
timestamp 1644511149
transform 1 0 29348 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_309
timestamp 1644511149
transform 1 0 29532 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_321
timestamp 1644511149
transform 1 0 30636 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_333
timestamp 1644511149
transform 1 0 31740 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_345
timestamp 1644511149
transform 1 0 32844 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_357
timestamp 1644511149
transform 1 0 33948 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_363
timestamp 1644511149
transform 1 0 34500 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_365
timestamp 1644511149
transform 1 0 34684 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_377
timestamp 1644511149
transform 1 0 35788 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_389
timestamp 1644511149
transform 1 0 36892 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_401
timestamp 1644511149
transform 1 0 37996 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_413
timestamp 1644511149
transform 1 0 39100 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_419
timestamp 1644511149
transform 1 0 39652 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_421
timestamp 1644511149
transform 1 0 39836 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_433
timestamp 1644511149
transform 1 0 40940 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_445
timestamp 1644511149
transform 1 0 42044 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_457
timestamp 1644511149
transform 1 0 43148 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_469
timestamp 1644511149
transform 1 0 44252 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_475
timestamp 1644511149
transform 1 0 44804 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_477
timestamp 1644511149
transform 1 0 44988 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_489
timestamp 1644511149
transform 1 0 46092 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_501
timestamp 1644511149
transform 1 0 47196 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_513
timestamp 1644511149
transform 1 0 48300 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_525
timestamp 1644511149
transform 1 0 49404 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_531
timestamp 1644511149
transform 1 0 49956 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_533
timestamp 1644511149
transform 1 0 50140 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_545
timestamp 1644511149
transform 1 0 51244 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_557
timestamp 1644511149
transform 1 0 52348 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_569
timestamp 1644511149
transform 1 0 53452 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_581
timestamp 1644511149
transform 1 0 54556 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_587
timestamp 1644511149
transform 1 0 55108 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_589
timestamp 1644511149
transform 1 0 55292 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_601
timestamp 1644511149
transform 1 0 56396 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_613
timestamp 1644511149
transform 1 0 57500 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_625
timestamp 1644511149
transform 1 0 58604 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_637
timestamp 1644511149
transform 1 0 59708 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_643
timestamp 1644511149
transform 1 0 60260 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_645
timestamp 1644511149
transform 1 0 60444 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_657
timestamp 1644511149
transform 1 0 61548 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_669
timestamp 1644511149
transform 1 0 62652 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_681
timestamp 1644511149
transform 1 0 63756 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_693
timestamp 1644511149
transform 1 0 64860 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_699
timestamp 1644511149
transform 1 0 65412 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_701
timestamp 1644511149
transform 1 0 65596 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_713
timestamp 1644511149
transform 1 0 66700 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_725
timestamp 1644511149
transform 1 0 67804 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_737
timestamp 1644511149
transform 1 0 68908 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_749
timestamp 1644511149
transform 1 0 70012 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_755
timestamp 1644511149
transform 1 0 70564 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_757
timestamp 1644511149
transform 1 0 70748 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_769
timestamp 1644511149
transform 1 0 71852 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_781
timestamp 1644511149
transform 1 0 72956 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_793
timestamp 1644511149
transform 1 0 74060 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_805
timestamp 1644511149
transform 1 0 75164 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_811
timestamp 1644511149
transform 1 0 75716 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_813
timestamp 1644511149
transform 1 0 75900 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_825
timestamp 1644511149
transform 1 0 77004 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_78_837
timestamp 1644511149
transform 1 0 78108 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_78_841
timestamp 1644511149
transform 1 0 78476 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_3
timestamp 1644511149
transform 1 0 1380 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_15
timestamp 1644511149
transform 1 0 2484 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_27
timestamp 1644511149
transform 1 0 3588 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_39
timestamp 1644511149
transform 1 0 4692 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_79_51
timestamp 1644511149
transform 1 0 5796 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_55
timestamp 1644511149
transform 1 0 6164 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_57
timestamp 1644511149
transform 1 0 6348 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_69
timestamp 1644511149
transform 1 0 7452 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_81
timestamp 1644511149
transform 1 0 8556 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_93
timestamp 1644511149
transform 1 0 9660 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_105
timestamp 1644511149
transform 1 0 10764 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_111
timestamp 1644511149
transform 1 0 11316 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_113
timestamp 1644511149
transform 1 0 11500 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_125
timestamp 1644511149
transform 1 0 12604 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_137
timestamp 1644511149
transform 1 0 13708 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_149
timestamp 1644511149
transform 1 0 14812 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_161
timestamp 1644511149
transform 1 0 15916 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_167
timestamp 1644511149
transform 1 0 16468 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_169
timestamp 1644511149
transform 1 0 16652 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_181
timestamp 1644511149
transform 1 0 17756 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_193
timestamp 1644511149
transform 1 0 18860 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_205
timestamp 1644511149
transform 1 0 19964 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_217
timestamp 1644511149
transform 1 0 21068 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_223
timestamp 1644511149
transform 1 0 21620 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_225
timestamp 1644511149
transform 1 0 21804 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_237
timestamp 1644511149
transform 1 0 22908 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_249
timestamp 1644511149
transform 1 0 24012 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_261
timestamp 1644511149
transform 1 0 25116 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_273
timestamp 1644511149
transform 1 0 26220 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_279
timestamp 1644511149
transform 1 0 26772 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_281
timestamp 1644511149
transform 1 0 26956 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_293
timestamp 1644511149
transform 1 0 28060 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_305
timestamp 1644511149
transform 1 0 29164 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_317
timestamp 1644511149
transform 1 0 30268 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_329
timestamp 1644511149
transform 1 0 31372 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_335
timestamp 1644511149
transform 1 0 31924 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_337
timestamp 1644511149
transform 1 0 32108 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_349
timestamp 1644511149
transform 1 0 33212 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_361
timestamp 1644511149
transform 1 0 34316 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_373
timestamp 1644511149
transform 1 0 35420 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_385
timestamp 1644511149
transform 1 0 36524 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_391
timestamp 1644511149
transform 1 0 37076 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_393
timestamp 1644511149
transform 1 0 37260 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_405
timestamp 1644511149
transform 1 0 38364 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_417
timestamp 1644511149
transform 1 0 39468 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_429
timestamp 1644511149
transform 1 0 40572 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_441
timestamp 1644511149
transform 1 0 41676 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_447
timestamp 1644511149
transform 1 0 42228 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_449
timestamp 1644511149
transform 1 0 42412 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_461
timestamp 1644511149
transform 1 0 43516 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_473
timestamp 1644511149
transform 1 0 44620 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_485
timestamp 1644511149
transform 1 0 45724 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_497
timestamp 1644511149
transform 1 0 46828 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_503
timestamp 1644511149
transform 1 0 47380 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_505
timestamp 1644511149
transform 1 0 47564 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_517
timestamp 1644511149
transform 1 0 48668 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_529
timestamp 1644511149
transform 1 0 49772 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_541
timestamp 1644511149
transform 1 0 50876 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_553
timestamp 1644511149
transform 1 0 51980 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_559
timestamp 1644511149
transform 1 0 52532 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_561
timestamp 1644511149
transform 1 0 52716 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_573
timestamp 1644511149
transform 1 0 53820 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_585
timestamp 1644511149
transform 1 0 54924 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_597
timestamp 1644511149
transform 1 0 56028 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_609
timestamp 1644511149
transform 1 0 57132 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_615
timestamp 1644511149
transform 1 0 57684 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_617
timestamp 1644511149
transform 1 0 57868 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_629
timestamp 1644511149
transform 1 0 58972 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_641
timestamp 1644511149
transform 1 0 60076 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_653
timestamp 1644511149
transform 1 0 61180 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_665
timestamp 1644511149
transform 1 0 62284 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_671
timestamp 1644511149
transform 1 0 62836 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_673
timestamp 1644511149
transform 1 0 63020 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_685
timestamp 1644511149
transform 1 0 64124 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_697
timestamp 1644511149
transform 1 0 65228 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_709
timestamp 1644511149
transform 1 0 66332 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_721
timestamp 1644511149
transform 1 0 67436 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_727
timestamp 1644511149
transform 1 0 67988 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_729
timestamp 1644511149
transform 1 0 68172 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_741
timestamp 1644511149
transform 1 0 69276 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_753
timestamp 1644511149
transform 1 0 70380 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_765
timestamp 1644511149
transform 1 0 71484 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_777
timestamp 1644511149
transform 1 0 72588 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_783
timestamp 1644511149
transform 1 0 73140 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_785
timestamp 1644511149
transform 1 0 73324 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_797
timestamp 1644511149
transform 1 0 74428 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_809
timestamp 1644511149
transform 1 0 75532 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_821
timestamp 1644511149
transform 1 0 76636 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_833
timestamp 1644511149
transform 1 0 77740 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_839
timestamp 1644511149
transform 1 0 78292 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_79_841
timestamp 1644511149
transform 1 0 78476 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_3
timestamp 1644511149
transform 1 0 1380 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_15
timestamp 1644511149
transform 1 0 2484 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_80_27
timestamp 1644511149
transform 1 0 3588 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_29
timestamp 1644511149
transform 1 0 3772 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_41
timestamp 1644511149
transform 1 0 4876 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_53
timestamp 1644511149
transform 1 0 5980 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_65
timestamp 1644511149
transform 1 0 7084 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_77
timestamp 1644511149
transform 1 0 8188 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_83
timestamp 1644511149
transform 1 0 8740 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_85
timestamp 1644511149
transform 1 0 8924 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_97
timestamp 1644511149
transform 1 0 10028 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_109
timestamp 1644511149
transform 1 0 11132 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_121
timestamp 1644511149
transform 1 0 12236 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_133
timestamp 1644511149
transform 1 0 13340 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_139
timestamp 1644511149
transform 1 0 13892 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_141
timestamp 1644511149
transform 1 0 14076 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_153
timestamp 1644511149
transform 1 0 15180 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_165
timestamp 1644511149
transform 1 0 16284 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_177
timestamp 1644511149
transform 1 0 17388 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_189
timestamp 1644511149
transform 1 0 18492 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_195
timestamp 1644511149
transform 1 0 19044 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_197
timestamp 1644511149
transform 1 0 19228 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_209
timestamp 1644511149
transform 1 0 20332 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_221
timestamp 1644511149
transform 1 0 21436 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_233
timestamp 1644511149
transform 1 0 22540 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_245
timestamp 1644511149
transform 1 0 23644 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_251
timestamp 1644511149
transform 1 0 24196 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_253
timestamp 1644511149
transform 1 0 24380 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_265
timestamp 1644511149
transform 1 0 25484 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_277
timestamp 1644511149
transform 1 0 26588 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_289
timestamp 1644511149
transform 1 0 27692 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_301
timestamp 1644511149
transform 1 0 28796 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_307
timestamp 1644511149
transform 1 0 29348 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_309
timestamp 1644511149
transform 1 0 29532 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_321
timestamp 1644511149
transform 1 0 30636 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_333
timestamp 1644511149
transform 1 0 31740 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_345
timestamp 1644511149
transform 1 0 32844 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_357
timestamp 1644511149
transform 1 0 33948 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_363
timestamp 1644511149
transform 1 0 34500 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_365
timestamp 1644511149
transform 1 0 34684 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_377
timestamp 1644511149
transform 1 0 35788 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_389
timestamp 1644511149
transform 1 0 36892 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_401
timestamp 1644511149
transform 1 0 37996 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_413
timestamp 1644511149
transform 1 0 39100 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_419
timestamp 1644511149
transform 1 0 39652 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_421
timestamp 1644511149
transform 1 0 39836 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_433
timestamp 1644511149
transform 1 0 40940 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_445
timestamp 1644511149
transform 1 0 42044 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_457
timestamp 1644511149
transform 1 0 43148 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_469
timestamp 1644511149
transform 1 0 44252 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_475
timestamp 1644511149
transform 1 0 44804 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_477
timestamp 1644511149
transform 1 0 44988 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_489
timestamp 1644511149
transform 1 0 46092 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_501
timestamp 1644511149
transform 1 0 47196 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_513
timestamp 1644511149
transform 1 0 48300 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_525
timestamp 1644511149
transform 1 0 49404 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_531
timestamp 1644511149
transform 1 0 49956 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_533
timestamp 1644511149
transform 1 0 50140 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_545
timestamp 1644511149
transform 1 0 51244 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_557
timestamp 1644511149
transform 1 0 52348 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_569
timestamp 1644511149
transform 1 0 53452 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_581
timestamp 1644511149
transform 1 0 54556 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_587
timestamp 1644511149
transform 1 0 55108 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_589
timestamp 1644511149
transform 1 0 55292 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_601
timestamp 1644511149
transform 1 0 56396 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_613
timestamp 1644511149
transform 1 0 57500 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_625
timestamp 1644511149
transform 1 0 58604 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_637
timestamp 1644511149
transform 1 0 59708 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_643
timestamp 1644511149
transform 1 0 60260 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_645
timestamp 1644511149
transform 1 0 60444 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_657
timestamp 1644511149
transform 1 0 61548 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_669
timestamp 1644511149
transform 1 0 62652 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_681
timestamp 1644511149
transform 1 0 63756 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_693
timestamp 1644511149
transform 1 0 64860 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_699
timestamp 1644511149
transform 1 0 65412 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_701
timestamp 1644511149
transform 1 0 65596 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_713
timestamp 1644511149
transform 1 0 66700 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_725
timestamp 1644511149
transform 1 0 67804 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_737
timestamp 1644511149
transform 1 0 68908 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_749
timestamp 1644511149
transform 1 0 70012 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_755
timestamp 1644511149
transform 1 0 70564 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_757
timestamp 1644511149
transform 1 0 70748 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_769
timestamp 1644511149
transform 1 0 71852 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_781
timestamp 1644511149
transform 1 0 72956 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_793
timestamp 1644511149
transform 1 0 74060 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_805
timestamp 1644511149
transform 1 0 75164 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_811
timestamp 1644511149
transform 1 0 75716 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_813
timestamp 1644511149
transform 1 0 75900 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_825
timestamp 1644511149
transform 1 0 77004 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_80_837
timestamp 1644511149
transform 1 0 78108 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_80_841
timestamp 1644511149
transform 1 0 78476 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_3
timestamp 1644511149
transform 1 0 1380 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_15
timestamp 1644511149
transform 1 0 2484 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_27
timestamp 1644511149
transform 1 0 3588 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_39
timestamp 1644511149
transform 1 0 4692 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_81_51
timestamp 1644511149
transform 1 0 5796 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_55
timestamp 1644511149
transform 1 0 6164 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_57
timestamp 1644511149
transform 1 0 6348 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_69
timestamp 1644511149
transform 1 0 7452 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_81
timestamp 1644511149
transform 1 0 8556 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_93
timestamp 1644511149
transform 1 0 9660 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_105
timestamp 1644511149
transform 1 0 10764 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_111
timestamp 1644511149
transform 1 0 11316 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_113
timestamp 1644511149
transform 1 0 11500 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_125
timestamp 1644511149
transform 1 0 12604 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_137
timestamp 1644511149
transform 1 0 13708 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_149
timestamp 1644511149
transform 1 0 14812 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_161
timestamp 1644511149
transform 1 0 15916 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_167
timestamp 1644511149
transform 1 0 16468 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_169
timestamp 1644511149
transform 1 0 16652 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_181
timestamp 1644511149
transform 1 0 17756 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_193
timestamp 1644511149
transform 1 0 18860 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_205
timestamp 1644511149
transform 1 0 19964 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_217
timestamp 1644511149
transform 1 0 21068 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_223
timestamp 1644511149
transform 1 0 21620 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_225
timestamp 1644511149
transform 1 0 21804 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_237
timestamp 1644511149
transform 1 0 22908 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_249
timestamp 1644511149
transform 1 0 24012 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_261
timestamp 1644511149
transform 1 0 25116 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_273
timestamp 1644511149
transform 1 0 26220 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_279
timestamp 1644511149
transform 1 0 26772 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_281
timestamp 1644511149
transform 1 0 26956 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_293
timestamp 1644511149
transform 1 0 28060 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_305
timestamp 1644511149
transform 1 0 29164 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_317
timestamp 1644511149
transform 1 0 30268 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_329
timestamp 1644511149
transform 1 0 31372 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_335
timestamp 1644511149
transform 1 0 31924 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_337
timestamp 1644511149
transform 1 0 32108 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_349
timestamp 1644511149
transform 1 0 33212 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_361
timestamp 1644511149
transform 1 0 34316 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_373
timestamp 1644511149
transform 1 0 35420 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_385
timestamp 1644511149
transform 1 0 36524 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_391
timestamp 1644511149
transform 1 0 37076 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_393
timestamp 1644511149
transform 1 0 37260 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_405
timestamp 1644511149
transform 1 0 38364 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_417
timestamp 1644511149
transform 1 0 39468 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_429
timestamp 1644511149
transform 1 0 40572 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_441
timestamp 1644511149
transform 1 0 41676 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_447
timestamp 1644511149
transform 1 0 42228 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_449
timestamp 1644511149
transform 1 0 42412 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_461
timestamp 1644511149
transform 1 0 43516 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_473
timestamp 1644511149
transform 1 0 44620 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_485
timestamp 1644511149
transform 1 0 45724 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_497
timestamp 1644511149
transform 1 0 46828 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_503
timestamp 1644511149
transform 1 0 47380 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_505
timestamp 1644511149
transform 1 0 47564 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_517
timestamp 1644511149
transform 1 0 48668 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_529
timestamp 1644511149
transform 1 0 49772 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_541
timestamp 1644511149
transform 1 0 50876 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_553
timestamp 1644511149
transform 1 0 51980 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_559
timestamp 1644511149
transform 1 0 52532 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_561
timestamp 1644511149
transform 1 0 52716 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_573
timestamp 1644511149
transform 1 0 53820 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_585
timestamp 1644511149
transform 1 0 54924 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_597
timestamp 1644511149
transform 1 0 56028 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_609
timestamp 1644511149
transform 1 0 57132 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_615
timestamp 1644511149
transform 1 0 57684 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_617
timestamp 1644511149
transform 1 0 57868 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_629
timestamp 1644511149
transform 1 0 58972 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_641
timestamp 1644511149
transform 1 0 60076 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_653
timestamp 1644511149
transform 1 0 61180 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_665
timestamp 1644511149
transform 1 0 62284 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_671
timestamp 1644511149
transform 1 0 62836 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_673
timestamp 1644511149
transform 1 0 63020 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_685
timestamp 1644511149
transform 1 0 64124 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_697
timestamp 1644511149
transform 1 0 65228 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_709
timestamp 1644511149
transform 1 0 66332 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_721
timestamp 1644511149
transform 1 0 67436 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_727
timestamp 1644511149
transform 1 0 67988 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_729
timestamp 1644511149
transform 1 0 68172 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_741
timestamp 1644511149
transform 1 0 69276 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_753
timestamp 1644511149
transform 1 0 70380 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_765
timestamp 1644511149
transform 1 0 71484 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_777
timestamp 1644511149
transform 1 0 72588 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_783
timestamp 1644511149
transform 1 0 73140 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_785
timestamp 1644511149
transform 1 0 73324 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_797
timestamp 1644511149
transform 1 0 74428 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_809
timestamp 1644511149
transform 1 0 75532 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_821
timestamp 1644511149
transform 1 0 76636 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_833
timestamp 1644511149
transform 1 0 77740 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_839
timestamp 1644511149
transform 1 0 78292 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_81_841
timestamp 1644511149
transform 1 0 78476 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_82_7
timestamp 1644511149
transform 1 0 1748 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_82_19
timestamp 1644511149
transform 1 0 2852 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_82_27
timestamp 1644511149
transform 1 0 3588 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_82_29
timestamp 1644511149
transform 1 0 3772 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_41
timestamp 1644511149
transform 1 0 4876 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_53
timestamp 1644511149
transform 1 0 5980 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_65
timestamp 1644511149
transform 1 0 7084 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_77
timestamp 1644511149
transform 1 0 8188 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_83
timestamp 1644511149
transform 1 0 8740 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_82_85
timestamp 1644511149
transform 1 0 8924 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_97
timestamp 1644511149
transform 1 0 10028 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_109
timestamp 1644511149
transform 1 0 11132 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_121
timestamp 1644511149
transform 1 0 12236 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_133
timestamp 1644511149
transform 1 0 13340 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_139
timestamp 1644511149
transform 1 0 13892 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_82_141
timestamp 1644511149
transform 1 0 14076 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_153
timestamp 1644511149
transform 1 0 15180 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_165
timestamp 1644511149
transform 1 0 16284 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_177
timestamp 1644511149
transform 1 0 17388 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_189
timestamp 1644511149
transform 1 0 18492 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_195
timestamp 1644511149
transform 1 0 19044 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_82_197
timestamp 1644511149
transform 1 0 19228 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_209
timestamp 1644511149
transform 1 0 20332 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_221
timestamp 1644511149
transform 1 0 21436 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_233
timestamp 1644511149
transform 1 0 22540 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_245
timestamp 1644511149
transform 1 0 23644 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_251
timestamp 1644511149
transform 1 0 24196 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_82_253
timestamp 1644511149
transform 1 0 24380 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_265
timestamp 1644511149
transform 1 0 25484 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_277
timestamp 1644511149
transform 1 0 26588 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_289
timestamp 1644511149
transform 1 0 27692 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_301
timestamp 1644511149
transform 1 0 28796 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_307
timestamp 1644511149
transform 1 0 29348 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_82_309
timestamp 1644511149
transform 1 0 29532 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_321
timestamp 1644511149
transform 1 0 30636 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_333
timestamp 1644511149
transform 1 0 31740 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_345
timestamp 1644511149
transform 1 0 32844 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_357
timestamp 1644511149
transform 1 0 33948 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_363
timestamp 1644511149
transform 1 0 34500 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_82_365
timestamp 1644511149
transform 1 0 34684 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_377
timestamp 1644511149
transform 1 0 35788 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_389
timestamp 1644511149
transform 1 0 36892 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_401
timestamp 1644511149
transform 1 0 37996 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_413
timestamp 1644511149
transform 1 0 39100 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_419
timestamp 1644511149
transform 1 0 39652 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_82_421
timestamp 1644511149
transform 1 0 39836 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_433
timestamp 1644511149
transform 1 0 40940 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_445
timestamp 1644511149
transform 1 0 42044 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_457
timestamp 1644511149
transform 1 0 43148 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_469
timestamp 1644511149
transform 1 0 44252 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_475
timestamp 1644511149
transform 1 0 44804 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_82_477
timestamp 1644511149
transform 1 0 44988 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_489
timestamp 1644511149
transform 1 0 46092 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_501
timestamp 1644511149
transform 1 0 47196 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_513
timestamp 1644511149
transform 1 0 48300 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_525
timestamp 1644511149
transform 1 0 49404 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_531
timestamp 1644511149
transform 1 0 49956 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_82_533
timestamp 1644511149
transform 1 0 50140 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_545
timestamp 1644511149
transform 1 0 51244 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_557
timestamp 1644511149
transform 1 0 52348 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_569
timestamp 1644511149
transform 1 0 53452 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_581
timestamp 1644511149
transform 1 0 54556 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_587
timestamp 1644511149
transform 1 0 55108 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_82_589
timestamp 1644511149
transform 1 0 55292 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_601
timestamp 1644511149
transform 1 0 56396 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_613
timestamp 1644511149
transform 1 0 57500 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_625
timestamp 1644511149
transform 1 0 58604 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_637
timestamp 1644511149
transform 1 0 59708 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_643
timestamp 1644511149
transform 1 0 60260 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_82_645
timestamp 1644511149
transform 1 0 60444 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_657
timestamp 1644511149
transform 1 0 61548 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_669
timestamp 1644511149
transform 1 0 62652 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_681
timestamp 1644511149
transform 1 0 63756 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_693
timestamp 1644511149
transform 1 0 64860 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_699
timestamp 1644511149
transform 1 0 65412 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_82_701
timestamp 1644511149
transform 1 0 65596 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_713
timestamp 1644511149
transform 1 0 66700 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_725
timestamp 1644511149
transform 1 0 67804 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_737
timestamp 1644511149
transform 1 0 68908 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_749
timestamp 1644511149
transform 1 0 70012 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_755
timestamp 1644511149
transform 1 0 70564 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_82_757
timestamp 1644511149
transform 1 0 70748 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_769
timestamp 1644511149
transform 1 0 71852 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_781
timestamp 1644511149
transform 1 0 72956 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_793
timestamp 1644511149
transform 1 0 74060 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_805
timestamp 1644511149
transform 1 0 75164 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_811
timestamp 1644511149
transform 1 0 75716 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_82_813
timestamp 1644511149
transform 1 0 75900 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_825
timestamp 1644511149
transform 1 0 77004 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_82_837
timestamp 1644511149
transform 1 0 78108 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_82_841
timestamp 1644511149
transform 1 0 78476 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_83_3
timestamp 1644511149
transform 1 0 1380 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_15
timestamp 1644511149
transform 1 0 2484 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_27
timestamp 1644511149
transform 1 0 3588 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_39
timestamp 1644511149
transform 1 0 4692 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_83_51
timestamp 1644511149
transform 1 0 5796 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_83_55
timestamp 1644511149
transform 1 0 6164 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_83_57
timestamp 1644511149
transform 1 0 6348 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_69
timestamp 1644511149
transform 1 0 7452 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_81
timestamp 1644511149
transform 1 0 8556 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_93
timestamp 1644511149
transform 1 0 9660 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_105
timestamp 1644511149
transform 1 0 10764 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_111
timestamp 1644511149
transform 1 0 11316 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_83_113
timestamp 1644511149
transform 1 0 11500 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_125
timestamp 1644511149
transform 1 0 12604 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_137
timestamp 1644511149
transform 1 0 13708 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_149
timestamp 1644511149
transform 1 0 14812 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_161
timestamp 1644511149
transform 1 0 15916 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_167
timestamp 1644511149
transform 1 0 16468 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_83_169
timestamp 1644511149
transform 1 0 16652 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_181
timestamp 1644511149
transform 1 0 17756 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_193
timestamp 1644511149
transform 1 0 18860 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_205
timestamp 1644511149
transform 1 0 19964 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_217
timestamp 1644511149
transform 1 0 21068 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_223
timestamp 1644511149
transform 1 0 21620 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_83_225
timestamp 1644511149
transform 1 0 21804 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_237
timestamp 1644511149
transform 1 0 22908 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_249
timestamp 1644511149
transform 1 0 24012 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_261
timestamp 1644511149
transform 1 0 25116 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_273
timestamp 1644511149
transform 1 0 26220 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_279
timestamp 1644511149
transform 1 0 26772 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_83_281
timestamp 1644511149
transform 1 0 26956 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_293
timestamp 1644511149
transform 1 0 28060 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_305
timestamp 1644511149
transform 1 0 29164 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_317
timestamp 1644511149
transform 1 0 30268 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_329
timestamp 1644511149
transform 1 0 31372 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_335
timestamp 1644511149
transform 1 0 31924 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_83_337
timestamp 1644511149
transform 1 0 32108 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_349
timestamp 1644511149
transform 1 0 33212 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_361
timestamp 1644511149
transform 1 0 34316 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_373
timestamp 1644511149
transform 1 0 35420 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_385
timestamp 1644511149
transform 1 0 36524 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_391
timestamp 1644511149
transform 1 0 37076 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_83_393
timestamp 1644511149
transform 1 0 37260 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_405
timestamp 1644511149
transform 1 0 38364 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_417
timestamp 1644511149
transform 1 0 39468 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_429
timestamp 1644511149
transform 1 0 40572 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_441
timestamp 1644511149
transform 1 0 41676 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_447
timestamp 1644511149
transform 1 0 42228 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_83_449
timestamp 1644511149
transform 1 0 42412 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_461
timestamp 1644511149
transform 1 0 43516 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_473
timestamp 1644511149
transform 1 0 44620 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_485
timestamp 1644511149
transform 1 0 45724 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_497
timestamp 1644511149
transform 1 0 46828 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_503
timestamp 1644511149
transform 1 0 47380 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_83_505
timestamp 1644511149
transform 1 0 47564 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_517
timestamp 1644511149
transform 1 0 48668 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_529
timestamp 1644511149
transform 1 0 49772 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_541
timestamp 1644511149
transform 1 0 50876 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_553
timestamp 1644511149
transform 1 0 51980 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_559
timestamp 1644511149
transform 1 0 52532 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_83_561
timestamp 1644511149
transform 1 0 52716 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_573
timestamp 1644511149
transform 1 0 53820 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_585
timestamp 1644511149
transform 1 0 54924 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_597
timestamp 1644511149
transform 1 0 56028 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_609
timestamp 1644511149
transform 1 0 57132 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_615
timestamp 1644511149
transform 1 0 57684 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_83_617
timestamp 1644511149
transform 1 0 57868 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_629
timestamp 1644511149
transform 1 0 58972 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_641
timestamp 1644511149
transform 1 0 60076 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_653
timestamp 1644511149
transform 1 0 61180 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_665
timestamp 1644511149
transform 1 0 62284 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_671
timestamp 1644511149
transform 1 0 62836 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_83_673
timestamp 1644511149
transform 1 0 63020 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_685
timestamp 1644511149
transform 1 0 64124 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_697
timestamp 1644511149
transform 1 0 65228 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_709
timestamp 1644511149
transform 1 0 66332 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_721
timestamp 1644511149
transform 1 0 67436 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_727
timestamp 1644511149
transform 1 0 67988 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_83_729
timestamp 1644511149
transform 1 0 68172 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_741
timestamp 1644511149
transform 1 0 69276 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_753
timestamp 1644511149
transform 1 0 70380 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_765
timestamp 1644511149
transform 1 0 71484 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_777
timestamp 1644511149
transform 1 0 72588 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_783
timestamp 1644511149
transform 1 0 73140 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_83_785
timestamp 1644511149
transform 1 0 73324 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_797
timestamp 1644511149
transform 1 0 74428 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_809
timestamp 1644511149
transform 1 0 75532 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_821
timestamp 1644511149
transform 1 0 76636 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_833
timestamp 1644511149
transform 1 0 77740 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_839
timestamp 1644511149
transform 1 0 78292 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_83_841
timestamp 1644511149
transform 1 0 78476 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_84_3
timestamp 1644511149
transform 1 0 1380 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_15
timestamp 1644511149
transform 1 0 2484 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_84_27
timestamp 1644511149
transform 1 0 3588 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_84_29
timestamp 1644511149
transform 1 0 3772 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_41
timestamp 1644511149
transform 1 0 4876 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_53
timestamp 1644511149
transform 1 0 5980 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_65
timestamp 1644511149
transform 1 0 7084 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_77
timestamp 1644511149
transform 1 0 8188 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_83
timestamp 1644511149
transform 1 0 8740 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_84_85
timestamp 1644511149
transform 1 0 8924 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_97
timestamp 1644511149
transform 1 0 10028 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_109
timestamp 1644511149
transform 1 0 11132 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_121
timestamp 1644511149
transform 1 0 12236 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_133
timestamp 1644511149
transform 1 0 13340 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_139
timestamp 1644511149
transform 1 0 13892 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_84_141
timestamp 1644511149
transform 1 0 14076 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_153
timestamp 1644511149
transform 1 0 15180 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_165
timestamp 1644511149
transform 1 0 16284 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_177
timestamp 1644511149
transform 1 0 17388 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_189
timestamp 1644511149
transform 1 0 18492 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_195
timestamp 1644511149
transform 1 0 19044 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_84_197
timestamp 1644511149
transform 1 0 19228 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_209
timestamp 1644511149
transform 1 0 20332 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_221
timestamp 1644511149
transform 1 0 21436 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_233
timestamp 1644511149
transform 1 0 22540 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_245
timestamp 1644511149
transform 1 0 23644 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_251
timestamp 1644511149
transform 1 0 24196 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_84_253
timestamp 1644511149
transform 1 0 24380 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_265
timestamp 1644511149
transform 1 0 25484 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_277
timestamp 1644511149
transform 1 0 26588 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_289
timestamp 1644511149
transform 1 0 27692 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_301
timestamp 1644511149
transform 1 0 28796 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_307
timestamp 1644511149
transform 1 0 29348 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_84_309
timestamp 1644511149
transform 1 0 29532 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_321
timestamp 1644511149
transform 1 0 30636 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_333
timestamp 1644511149
transform 1 0 31740 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_345
timestamp 1644511149
transform 1 0 32844 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_357
timestamp 1644511149
transform 1 0 33948 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_363
timestamp 1644511149
transform 1 0 34500 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_84_365
timestamp 1644511149
transform 1 0 34684 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_377
timestamp 1644511149
transform 1 0 35788 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_389
timestamp 1644511149
transform 1 0 36892 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_401
timestamp 1644511149
transform 1 0 37996 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_413
timestamp 1644511149
transform 1 0 39100 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_419
timestamp 1644511149
transform 1 0 39652 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_84_421
timestamp 1644511149
transform 1 0 39836 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_433
timestamp 1644511149
transform 1 0 40940 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_445
timestamp 1644511149
transform 1 0 42044 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_457
timestamp 1644511149
transform 1 0 43148 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_469
timestamp 1644511149
transform 1 0 44252 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_475
timestamp 1644511149
transform 1 0 44804 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_84_477
timestamp 1644511149
transform 1 0 44988 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_489
timestamp 1644511149
transform 1 0 46092 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_501
timestamp 1644511149
transform 1 0 47196 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_513
timestamp 1644511149
transform 1 0 48300 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_525
timestamp 1644511149
transform 1 0 49404 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_531
timestamp 1644511149
transform 1 0 49956 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_84_533
timestamp 1644511149
transform 1 0 50140 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_545
timestamp 1644511149
transform 1 0 51244 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_557
timestamp 1644511149
transform 1 0 52348 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_569
timestamp 1644511149
transform 1 0 53452 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_581
timestamp 1644511149
transform 1 0 54556 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_587
timestamp 1644511149
transform 1 0 55108 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_84_589
timestamp 1644511149
transform 1 0 55292 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_601
timestamp 1644511149
transform 1 0 56396 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_613
timestamp 1644511149
transform 1 0 57500 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_625
timestamp 1644511149
transform 1 0 58604 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_637
timestamp 1644511149
transform 1 0 59708 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_643
timestamp 1644511149
transform 1 0 60260 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_84_645
timestamp 1644511149
transform 1 0 60444 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_657
timestamp 1644511149
transform 1 0 61548 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_669
timestamp 1644511149
transform 1 0 62652 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_681
timestamp 1644511149
transform 1 0 63756 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_693
timestamp 1644511149
transform 1 0 64860 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_699
timestamp 1644511149
transform 1 0 65412 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_84_701
timestamp 1644511149
transform 1 0 65596 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_713
timestamp 1644511149
transform 1 0 66700 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_725
timestamp 1644511149
transform 1 0 67804 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_737
timestamp 1644511149
transform 1 0 68908 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_749
timestamp 1644511149
transform 1 0 70012 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_755
timestamp 1644511149
transform 1 0 70564 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_84_757
timestamp 1644511149
transform 1 0 70748 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_769
timestamp 1644511149
transform 1 0 71852 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_781
timestamp 1644511149
transform 1 0 72956 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_793
timestamp 1644511149
transform 1 0 74060 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_805
timestamp 1644511149
transform 1 0 75164 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_811
timestamp 1644511149
transform 1 0 75716 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_84_813
timestamp 1644511149
transform 1 0 75900 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_825
timestamp 1644511149
transform 1 0 77004 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_84_837
timestamp 1644511149
transform 1 0 78108 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_84_841
timestamp 1644511149
transform 1 0 78476 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_85_3
timestamp 1644511149
transform 1 0 1380 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_15
timestamp 1644511149
transform 1 0 2484 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_27
timestamp 1644511149
transform 1 0 3588 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_39
timestamp 1644511149
transform 1 0 4692 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_85_51
timestamp 1644511149
transform 1 0 5796 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_85_55
timestamp 1644511149
transform 1 0 6164 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_85_57
timestamp 1644511149
transform 1 0 6348 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_69
timestamp 1644511149
transform 1 0 7452 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_81
timestamp 1644511149
transform 1 0 8556 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_93
timestamp 1644511149
transform 1 0 9660 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_105
timestamp 1644511149
transform 1 0 10764 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_111
timestamp 1644511149
transform 1 0 11316 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_85_113
timestamp 1644511149
transform 1 0 11500 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_125
timestamp 1644511149
transform 1 0 12604 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_137
timestamp 1644511149
transform 1 0 13708 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_149
timestamp 1644511149
transform 1 0 14812 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_161
timestamp 1644511149
transform 1 0 15916 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_167
timestamp 1644511149
transform 1 0 16468 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_85_169
timestamp 1644511149
transform 1 0 16652 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_181
timestamp 1644511149
transform 1 0 17756 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_193
timestamp 1644511149
transform 1 0 18860 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_205
timestamp 1644511149
transform 1 0 19964 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_217
timestamp 1644511149
transform 1 0 21068 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_223
timestamp 1644511149
transform 1 0 21620 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_85_225
timestamp 1644511149
transform 1 0 21804 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_237
timestamp 1644511149
transform 1 0 22908 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_249
timestamp 1644511149
transform 1 0 24012 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_261
timestamp 1644511149
transform 1 0 25116 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_273
timestamp 1644511149
transform 1 0 26220 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_279
timestamp 1644511149
transform 1 0 26772 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_85_281
timestamp 1644511149
transform 1 0 26956 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_293
timestamp 1644511149
transform 1 0 28060 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_305
timestamp 1644511149
transform 1 0 29164 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_317
timestamp 1644511149
transform 1 0 30268 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_329
timestamp 1644511149
transform 1 0 31372 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_335
timestamp 1644511149
transform 1 0 31924 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_85_337
timestamp 1644511149
transform 1 0 32108 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_349
timestamp 1644511149
transform 1 0 33212 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_361
timestamp 1644511149
transform 1 0 34316 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_373
timestamp 1644511149
transform 1 0 35420 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_385
timestamp 1644511149
transform 1 0 36524 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_391
timestamp 1644511149
transform 1 0 37076 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_85_393
timestamp 1644511149
transform 1 0 37260 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_405
timestamp 1644511149
transform 1 0 38364 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_417
timestamp 1644511149
transform 1 0 39468 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_429
timestamp 1644511149
transform 1 0 40572 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_441
timestamp 1644511149
transform 1 0 41676 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_447
timestamp 1644511149
transform 1 0 42228 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_85_449
timestamp 1644511149
transform 1 0 42412 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_461
timestamp 1644511149
transform 1 0 43516 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_473
timestamp 1644511149
transform 1 0 44620 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_485
timestamp 1644511149
transform 1 0 45724 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_497
timestamp 1644511149
transform 1 0 46828 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_503
timestamp 1644511149
transform 1 0 47380 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_85_505
timestamp 1644511149
transform 1 0 47564 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_517
timestamp 1644511149
transform 1 0 48668 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_529
timestamp 1644511149
transform 1 0 49772 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_541
timestamp 1644511149
transform 1 0 50876 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_553
timestamp 1644511149
transform 1 0 51980 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_559
timestamp 1644511149
transform 1 0 52532 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_85_561
timestamp 1644511149
transform 1 0 52716 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_573
timestamp 1644511149
transform 1 0 53820 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_585
timestamp 1644511149
transform 1 0 54924 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_597
timestamp 1644511149
transform 1 0 56028 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_609
timestamp 1644511149
transform 1 0 57132 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_615
timestamp 1644511149
transform 1 0 57684 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_85_617
timestamp 1644511149
transform 1 0 57868 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_629
timestamp 1644511149
transform 1 0 58972 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_641
timestamp 1644511149
transform 1 0 60076 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_653
timestamp 1644511149
transform 1 0 61180 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_665
timestamp 1644511149
transform 1 0 62284 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_671
timestamp 1644511149
transform 1 0 62836 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_85_673
timestamp 1644511149
transform 1 0 63020 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_685
timestamp 1644511149
transform 1 0 64124 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_697
timestamp 1644511149
transform 1 0 65228 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_709
timestamp 1644511149
transform 1 0 66332 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_721
timestamp 1644511149
transform 1 0 67436 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_727
timestamp 1644511149
transform 1 0 67988 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_85_729
timestamp 1644511149
transform 1 0 68172 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_741
timestamp 1644511149
transform 1 0 69276 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_753
timestamp 1644511149
transform 1 0 70380 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_765
timestamp 1644511149
transform 1 0 71484 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_777
timestamp 1644511149
transform 1 0 72588 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_783
timestamp 1644511149
transform 1 0 73140 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_85_785
timestamp 1644511149
transform 1 0 73324 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_797
timestamp 1644511149
transform 1 0 74428 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_809
timestamp 1644511149
transform 1 0 75532 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_821
timestamp 1644511149
transform 1 0 76636 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_833
timestamp 1644511149
transform 1 0 77740 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_839
timestamp 1644511149
transform 1 0 78292 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_85_841
timestamp 1644511149
transform 1 0 78476 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_86_3
timestamp 1644511149
transform 1 0 1380 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_15
timestamp 1644511149
transform 1 0 2484 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_86_27
timestamp 1644511149
transform 1 0 3588 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_86_29
timestamp 1644511149
transform 1 0 3772 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_41
timestamp 1644511149
transform 1 0 4876 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_53
timestamp 1644511149
transform 1 0 5980 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_65
timestamp 1644511149
transform 1 0 7084 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_77
timestamp 1644511149
transform 1 0 8188 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_83
timestamp 1644511149
transform 1 0 8740 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_86_85
timestamp 1644511149
transform 1 0 8924 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_97
timestamp 1644511149
transform 1 0 10028 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_109
timestamp 1644511149
transform 1 0 11132 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_121
timestamp 1644511149
transform 1 0 12236 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_133
timestamp 1644511149
transform 1 0 13340 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_139
timestamp 1644511149
transform 1 0 13892 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_86_141
timestamp 1644511149
transform 1 0 14076 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_153
timestamp 1644511149
transform 1 0 15180 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_165
timestamp 1644511149
transform 1 0 16284 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_177
timestamp 1644511149
transform 1 0 17388 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_189
timestamp 1644511149
transform 1 0 18492 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_195
timestamp 1644511149
transform 1 0 19044 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_86_197
timestamp 1644511149
transform 1 0 19228 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_209
timestamp 1644511149
transform 1 0 20332 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_221
timestamp 1644511149
transform 1 0 21436 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_233
timestamp 1644511149
transform 1 0 22540 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_245
timestamp 1644511149
transform 1 0 23644 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_251
timestamp 1644511149
transform 1 0 24196 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_86_253
timestamp 1644511149
transform 1 0 24380 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_265
timestamp 1644511149
transform 1 0 25484 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_277
timestamp 1644511149
transform 1 0 26588 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_289
timestamp 1644511149
transform 1 0 27692 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_301
timestamp 1644511149
transform 1 0 28796 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_307
timestamp 1644511149
transform 1 0 29348 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_86_309
timestamp 1644511149
transform 1 0 29532 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_321
timestamp 1644511149
transform 1 0 30636 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_333
timestamp 1644511149
transform 1 0 31740 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_345
timestamp 1644511149
transform 1 0 32844 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_357
timestamp 1644511149
transform 1 0 33948 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_363
timestamp 1644511149
transform 1 0 34500 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_86_365
timestamp 1644511149
transform 1 0 34684 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_377
timestamp 1644511149
transform 1 0 35788 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_389
timestamp 1644511149
transform 1 0 36892 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_401
timestamp 1644511149
transform 1 0 37996 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_413
timestamp 1644511149
transform 1 0 39100 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_419
timestamp 1644511149
transform 1 0 39652 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_86_421
timestamp 1644511149
transform 1 0 39836 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_433
timestamp 1644511149
transform 1 0 40940 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_445
timestamp 1644511149
transform 1 0 42044 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_457
timestamp 1644511149
transform 1 0 43148 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_469
timestamp 1644511149
transform 1 0 44252 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_475
timestamp 1644511149
transform 1 0 44804 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_86_477
timestamp 1644511149
transform 1 0 44988 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_489
timestamp 1644511149
transform 1 0 46092 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_501
timestamp 1644511149
transform 1 0 47196 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_513
timestamp 1644511149
transform 1 0 48300 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_525
timestamp 1644511149
transform 1 0 49404 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_531
timestamp 1644511149
transform 1 0 49956 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_86_533
timestamp 1644511149
transform 1 0 50140 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_545
timestamp 1644511149
transform 1 0 51244 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_557
timestamp 1644511149
transform 1 0 52348 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_569
timestamp 1644511149
transform 1 0 53452 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_581
timestamp 1644511149
transform 1 0 54556 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_587
timestamp 1644511149
transform 1 0 55108 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_86_589
timestamp 1644511149
transform 1 0 55292 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_601
timestamp 1644511149
transform 1 0 56396 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_613
timestamp 1644511149
transform 1 0 57500 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_625
timestamp 1644511149
transform 1 0 58604 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_637
timestamp 1644511149
transform 1 0 59708 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_643
timestamp 1644511149
transform 1 0 60260 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_86_645
timestamp 1644511149
transform 1 0 60444 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_657
timestamp 1644511149
transform 1 0 61548 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_669
timestamp 1644511149
transform 1 0 62652 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_681
timestamp 1644511149
transform 1 0 63756 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_693
timestamp 1644511149
transform 1 0 64860 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_699
timestamp 1644511149
transform 1 0 65412 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_86_701
timestamp 1644511149
transform 1 0 65596 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_713
timestamp 1644511149
transform 1 0 66700 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_725
timestamp 1644511149
transform 1 0 67804 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_737
timestamp 1644511149
transform 1 0 68908 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_749
timestamp 1644511149
transform 1 0 70012 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_755
timestamp 1644511149
transform 1 0 70564 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_86_757
timestamp 1644511149
transform 1 0 70748 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_769
timestamp 1644511149
transform 1 0 71852 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_781
timestamp 1644511149
transform 1 0 72956 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_793
timestamp 1644511149
transform 1 0 74060 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_805
timestamp 1644511149
transform 1 0 75164 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_811
timestamp 1644511149
transform 1 0 75716 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_86_813
timestamp 1644511149
transform 1 0 75900 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_825
timestamp 1644511149
transform 1 0 77004 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_86_837
timestamp 1644511149
transform 1 0 78108 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_86_841
timestamp 1644511149
transform 1 0 78476 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_87_3
timestamp 1644511149
transform 1 0 1380 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_15
timestamp 1644511149
transform 1 0 2484 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_27
timestamp 1644511149
transform 1 0 3588 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_39
timestamp 1644511149
transform 1 0 4692 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_87_51
timestamp 1644511149
transform 1 0 5796 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_87_55
timestamp 1644511149
transform 1 0 6164 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_87_57
timestamp 1644511149
transform 1 0 6348 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_69
timestamp 1644511149
transform 1 0 7452 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_81
timestamp 1644511149
transform 1 0 8556 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_93
timestamp 1644511149
transform 1 0 9660 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_105
timestamp 1644511149
transform 1 0 10764 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_111
timestamp 1644511149
transform 1 0 11316 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_87_113
timestamp 1644511149
transform 1 0 11500 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_125
timestamp 1644511149
transform 1 0 12604 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_137
timestamp 1644511149
transform 1 0 13708 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_149
timestamp 1644511149
transform 1 0 14812 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_161
timestamp 1644511149
transform 1 0 15916 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_167
timestamp 1644511149
transform 1 0 16468 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_87_169
timestamp 1644511149
transform 1 0 16652 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_181
timestamp 1644511149
transform 1 0 17756 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_193
timestamp 1644511149
transform 1 0 18860 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_205
timestamp 1644511149
transform 1 0 19964 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_217
timestamp 1644511149
transform 1 0 21068 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_223
timestamp 1644511149
transform 1 0 21620 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_87_225
timestamp 1644511149
transform 1 0 21804 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_237
timestamp 1644511149
transform 1 0 22908 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_249
timestamp 1644511149
transform 1 0 24012 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_261
timestamp 1644511149
transform 1 0 25116 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_273
timestamp 1644511149
transform 1 0 26220 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_279
timestamp 1644511149
transform 1 0 26772 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_87_281
timestamp 1644511149
transform 1 0 26956 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_293
timestamp 1644511149
transform 1 0 28060 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_305
timestamp 1644511149
transform 1 0 29164 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_317
timestamp 1644511149
transform 1 0 30268 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_329
timestamp 1644511149
transform 1 0 31372 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_335
timestamp 1644511149
transform 1 0 31924 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_87_337
timestamp 1644511149
transform 1 0 32108 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_349
timestamp 1644511149
transform 1 0 33212 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_361
timestamp 1644511149
transform 1 0 34316 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_373
timestamp 1644511149
transform 1 0 35420 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_385
timestamp 1644511149
transform 1 0 36524 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_391
timestamp 1644511149
transform 1 0 37076 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_87_393
timestamp 1644511149
transform 1 0 37260 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_405
timestamp 1644511149
transform 1 0 38364 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_417
timestamp 1644511149
transform 1 0 39468 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_429
timestamp 1644511149
transform 1 0 40572 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_441
timestamp 1644511149
transform 1 0 41676 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_447
timestamp 1644511149
transform 1 0 42228 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_87_449
timestamp 1644511149
transform 1 0 42412 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_461
timestamp 1644511149
transform 1 0 43516 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_473
timestamp 1644511149
transform 1 0 44620 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_485
timestamp 1644511149
transform 1 0 45724 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_497
timestamp 1644511149
transform 1 0 46828 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_503
timestamp 1644511149
transform 1 0 47380 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_87_505
timestamp 1644511149
transform 1 0 47564 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_517
timestamp 1644511149
transform 1 0 48668 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_529
timestamp 1644511149
transform 1 0 49772 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_541
timestamp 1644511149
transform 1 0 50876 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_553
timestamp 1644511149
transform 1 0 51980 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_559
timestamp 1644511149
transform 1 0 52532 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_87_561
timestamp 1644511149
transform 1 0 52716 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_573
timestamp 1644511149
transform 1 0 53820 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_585
timestamp 1644511149
transform 1 0 54924 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_597
timestamp 1644511149
transform 1 0 56028 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_609
timestamp 1644511149
transform 1 0 57132 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_615
timestamp 1644511149
transform 1 0 57684 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_87_617
timestamp 1644511149
transform 1 0 57868 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_629
timestamp 1644511149
transform 1 0 58972 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_641
timestamp 1644511149
transform 1 0 60076 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_653
timestamp 1644511149
transform 1 0 61180 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_665
timestamp 1644511149
transform 1 0 62284 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_671
timestamp 1644511149
transform 1 0 62836 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_87_673
timestamp 1644511149
transform 1 0 63020 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_685
timestamp 1644511149
transform 1 0 64124 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_697
timestamp 1644511149
transform 1 0 65228 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_709
timestamp 1644511149
transform 1 0 66332 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_721
timestamp 1644511149
transform 1 0 67436 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_727
timestamp 1644511149
transform 1 0 67988 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_87_729
timestamp 1644511149
transform 1 0 68172 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_741
timestamp 1644511149
transform 1 0 69276 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_753
timestamp 1644511149
transform 1 0 70380 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_765
timestamp 1644511149
transform 1 0 71484 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_777
timestamp 1644511149
transform 1 0 72588 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_783
timestamp 1644511149
transform 1 0 73140 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_87_785
timestamp 1644511149
transform 1 0 73324 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_797
timestamp 1644511149
transform 1 0 74428 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_809
timestamp 1644511149
transform 1 0 75532 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_821
timestamp 1644511149
transform 1 0 76636 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_833
timestamp 1644511149
transform 1 0 77740 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_839
timestamp 1644511149
transform 1 0 78292 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_87_841
timestamp 1644511149
transform 1 0 78476 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_88_3
timestamp 1644511149
transform 1 0 1380 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_15
timestamp 1644511149
transform 1 0 2484 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_88_27
timestamp 1644511149
transform 1 0 3588 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_88_29
timestamp 1644511149
transform 1 0 3772 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_41
timestamp 1644511149
transform 1 0 4876 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_53
timestamp 1644511149
transform 1 0 5980 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_65
timestamp 1644511149
transform 1 0 7084 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_77
timestamp 1644511149
transform 1 0 8188 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_83
timestamp 1644511149
transform 1 0 8740 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_88_85
timestamp 1644511149
transform 1 0 8924 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_97
timestamp 1644511149
transform 1 0 10028 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_109
timestamp 1644511149
transform 1 0 11132 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_121
timestamp 1644511149
transform 1 0 12236 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_133
timestamp 1644511149
transform 1 0 13340 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_139
timestamp 1644511149
transform 1 0 13892 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_88_141
timestamp 1644511149
transform 1 0 14076 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_153
timestamp 1644511149
transform 1 0 15180 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_165
timestamp 1644511149
transform 1 0 16284 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_177
timestamp 1644511149
transform 1 0 17388 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_189
timestamp 1644511149
transform 1 0 18492 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_195
timestamp 1644511149
transform 1 0 19044 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_88_197
timestamp 1644511149
transform 1 0 19228 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_209
timestamp 1644511149
transform 1 0 20332 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_221
timestamp 1644511149
transform 1 0 21436 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_233
timestamp 1644511149
transform 1 0 22540 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_245
timestamp 1644511149
transform 1 0 23644 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_251
timestamp 1644511149
transform 1 0 24196 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_88_253
timestamp 1644511149
transform 1 0 24380 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_265
timestamp 1644511149
transform 1 0 25484 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_277
timestamp 1644511149
transform 1 0 26588 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_289
timestamp 1644511149
transform 1 0 27692 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_301
timestamp 1644511149
transform 1 0 28796 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_307
timestamp 1644511149
transform 1 0 29348 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_88_309
timestamp 1644511149
transform 1 0 29532 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_321
timestamp 1644511149
transform 1 0 30636 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_333
timestamp 1644511149
transform 1 0 31740 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_345
timestamp 1644511149
transform 1 0 32844 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_357
timestamp 1644511149
transform 1 0 33948 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_363
timestamp 1644511149
transform 1 0 34500 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_88_365
timestamp 1644511149
transform 1 0 34684 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_377
timestamp 1644511149
transform 1 0 35788 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_389
timestamp 1644511149
transform 1 0 36892 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_401
timestamp 1644511149
transform 1 0 37996 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_413
timestamp 1644511149
transform 1 0 39100 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_419
timestamp 1644511149
transform 1 0 39652 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_88_421
timestamp 1644511149
transform 1 0 39836 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_433
timestamp 1644511149
transform 1 0 40940 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_445
timestamp 1644511149
transform 1 0 42044 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_457
timestamp 1644511149
transform 1 0 43148 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_469
timestamp 1644511149
transform 1 0 44252 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_475
timestamp 1644511149
transform 1 0 44804 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_88_477
timestamp 1644511149
transform 1 0 44988 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_489
timestamp 1644511149
transform 1 0 46092 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_501
timestamp 1644511149
transform 1 0 47196 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_513
timestamp 1644511149
transform 1 0 48300 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_525
timestamp 1644511149
transform 1 0 49404 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_531
timestamp 1644511149
transform 1 0 49956 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_88_533
timestamp 1644511149
transform 1 0 50140 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_545
timestamp 1644511149
transform 1 0 51244 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_557
timestamp 1644511149
transform 1 0 52348 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_569
timestamp 1644511149
transform 1 0 53452 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_581
timestamp 1644511149
transform 1 0 54556 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_587
timestamp 1644511149
transform 1 0 55108 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_88_589
timestamp 1644511149
transform 1 0 55292 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_601
timestamp 1644511149
transform 1 0 56396 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_613
timestamp 1644511149
transform 1 0 57500 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_625
timestamp 1644511149
transform 1 0 58604 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_637
timestamp 1644511149
transform 1 0 59708 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_643
timestamp 1644511149
transform 1 0 60260 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_88_645
timestamp 1644511149
transform 1 0 60444 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_657
timestamp 1644511149
transform 1 0 61548 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_669
timestamp 1644511149
transform 1 0 62652 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_681
timestamp 1644511149
transform 1 0 63756 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_693
timestamp 1644511149
transform 1 0 64860 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_699
timestamp 1644511149
transform 1 0 65412 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_88_701
timestamp 1644511149
transform 1 0 65596 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_713
timestamp 1644511149
transform 1 0 66700 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_725
timestamp 1644511149
transform 1 0 67804 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_737
timestamp 1644511149
transform 1 0 68908 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_749
timestamp 1644511149
transform 1 0 70012 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_755
timestamp 1644511149
transform 1 0 70564 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_88_757
timestamp 1644511149
transform 1 0 70748 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_769
timestamp 1644511149
transform 1 0 71852 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_781
timestamp 1644511149
transform 1 0 72956 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_793
timestamp 1644511149
transform 1 0 74060 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_805
timestamp 1644511149
transform 1 0 75164 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_811
timestamp 1644511149
transform 1 0 75716 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_88_813
timestamp 1644511149
transform 1 0 75900 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_825
timestamp 1644511149
transform 1 0 77004 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_88_837
timestamp 1644511149
transform 1 0 78108 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_88_841
timestamp 1644511149
transform 1 0 78476 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_89_7
timestamp 1644511149
transform 1 0 1748 0 -1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_89_11
timestamp 1644511149
transform 1 0 2116 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_23
timestamp 1644511149
transform 1 0 3220 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_35
timestamp 1644511149
transform 1 0 4324 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_89_47
timestamp 1644511149
transform 1 0 5428 0 -1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_89_55
timestamp 1644511149
transform 1 0 6164 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_89_57
timestamp 1644511149
transform 1 0 6348 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_69
timestamp 1644511149
transform 1 0 7452 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_81
timestamp 1644511149
transform 1 0 8556 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_93
timestamp 1644511149
transform 1 0 9660 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_105
timestamp 1644511149
transform 1 0 10764 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_111
timestamp 1644511149
transform 1 0 11316 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_89_113
timestamp 1644511149
transform 1 0 11500 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_125
timestamp 1644511149
transform 1 0 12604 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_137
timestamp 1644511149
transform 1 0 13708 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_149
timestamp 1644511149
transform 1 0 14812 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_161
timestamp 1644511149
transform 1 0 15916 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_167
timestamp 1644511149
transform 1 0 16468 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_89_169
timestamp 1644511149
transform 1 0 16652 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_181
timestamp 1644511149
transform 1 0 17756 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_193
timestamp 1644511149
transform 1 0 18860 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_205
timestamp 1644511149
transform 1 0 19964 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_217
timestamp 1644511149
transform 1 0 21068 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_223
timestamp 1644511149
transform 1 0 21620 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_89_225
timestamp 1644511149
transform 1 0 21804 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_237
timestamp 1644511149
transform 1 0 22908 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_249
timestamp 1644511149
transform 1 0 24012 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_261
timestamp 1644511149
transform 1 0 25116 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_273
timestamp 1644511149
transform 1 0 26220 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_279
timestamp 1644511149
transform 1 0 26772 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_89_281
timestamp 1644511149
transform 1 0 26956 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_293
timestamp 1644511149
transform 1 0 28060 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_305
timestamp 1644511149
transform 1 0 29164 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_317
timestamp 1644511149
transform 1 0 30268 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_329
timestamp 1644511149
transform 1 0 31372 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_335
timestamp 1644511149
transform 1 0 31924 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_89_337
timestamp 1644511149
transform 1 0 32108 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_349
timestamp 1644511149
transform 1 0 33212 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_361
timestamp 1644511149
transform 1 0 34316 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_373
timestamp 1644511149
transform 1 0 35420 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_385
timestamp 1644511149
transform 1 0 36524 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_391
timestamp 1644511149
transform 1 0 37076 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_89_393
timestamp 1644511149
transform 1 0 37260 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_405
timestamp 1644511149
transform 1 0 38364 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_417
timestamp 1644511149
transform 1 0 39468 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_429
timestamp 1644511149
transform 1 0 40572 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_441
timestamp 1644511149
transform 1 0 41676 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_447
timestamp 1644511149
transform 1 0 42228 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_89_449
timestamp 1644511149
transform 1 0 42412 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_461
timestamp 1644511149
transform 1 0 43516 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_473
timestamp 1644511149
transform 1 0 44620 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_485
timestamp 1644511149
transform 1 0 45724 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_497
timestamp 1644511149
transform 1 0 46828 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_503
timestamp 1644511149
transform 1 0 47380 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_89_505
timestamp 1644511149
transform 1 0 47564 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_517
timestamp 1644511149
transform 1 0 48668 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_529
timestamp 1644511149
transform 1 0 49772 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_541
timestamp 1644511149
transform 1 0 50876 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_553
timestamp 1644511149
transform 1 0 51980 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_559
timestamp 1644511149
transform 1 0 52532 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_89_561
timestamp 1644511149
transform 1 0 52716 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_573
timestamp 1644511149
transform 1 0 53820 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_585
timestamp 1644511149
transform 1 0 54924 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_597
timestamp 1644511149
transform 1 0 56028 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_609
timestamp 1644511149
transform 1 0 57132 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_615
timestamp 1644511149
transform 1 0 57684 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_89_617
timestamp 1644511149
transform 1 0 57868 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_629
timestamp 1644511149
transform 1 0 58972 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_641
timestamp 1644511149
transform 1 0 60076 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_653
timestamp 1644511149
transform 1 0 61180 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_665
timestamp 1644511149
transform 1 0 62284 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_671
timestamp 1644511149
transform 1 0 62836 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_89_673
timestamp 1644511149
transform 1 0 63020 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_685
timestamp 1644511149
transform 1 0 64124 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_697
timestamp 1644511149
transform 1 0 65228 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_709
timestamp 1644511149
transform 1 0 66332 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_721
timestamp 1644511149
transform 1 0 67436 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_727
timestamp 1644511149
transform 1 0 67988 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_89_729
timestamp 1644511149
transform 1 0 68172 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_741
timestamp 1644511149
transform 1 0 69276 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_753
timestamp 1644511149
transform 1 0 70380 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_765
timestamp 1644511149
transform 1 0 71484 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_777
timestamp 1644511149
transform 1 0 72588 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_783
timestamp 1644511149
transform 1 0 73140 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_89_785
timestamp 1644511149
transform 1 0 73324 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_797
timestamp 1644511149
transform 1 0 74428 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_809
timestamp 1644511149
transform 1 0 75532 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_821
timestamp 1644511149
transform 1 0 76636 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_833
timestamp 1644511149
transform 1 0 77740 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_839
timestamp 1644511149
transform 1 0 78292 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_89_841
timestamp 1644511149
transform 1 0 78476 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_90_3
timestamp 1644511149
transform 1 0 1380 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_15
timestamp 1644511149
transform 1 0 2484 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_90_27
timestamp 1644511149
transform 1 0 3588 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_90_29
timestamp 1644511149
transform 1 0 3772 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_41
timestamp 1644511149
transform 1 0 4876 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_53
timestamp 1644511149
transform 1 0 5980 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_65
timestamp 1644511149
transform 1 0 7084 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_77
timestamp 1644511149
transform 1 0 8188 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_83
timestamp 1644511149
transform 1 0 8740 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_90_85
timestamp 1644511149
transform 1 0 8924 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_97
timestamp 1644511149
transform 1 0 10028 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_109
timestamp 1644511149
transform 1 0 11132 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_121
timestamp 1644511149
transform 1 0 12236 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_133
timestamp 1644511149
transform 1 0 13340 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_139
timestamp 1644511149
transform 1 0 13892 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_90_141
timestamp 1644511149
transform 1 0 14076 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_153
timestamp 1644511149
transform 1 0 15180 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_165
timestamp 1644511149
transform 1 0 16284 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_177
timestamp 1644511149
transform 1 0 17388 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_189
timestamp 1644511149
transform 1 0 18492 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_195
timestamp 1644511149
transform 1 0 19044 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_90_197
timestamp 1644511149
transform 1 0 19228 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_209
timestamp 1644511149
transform 1 0 20332 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_221
timestamp 1644511149
transform 1 0 21436 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_233
timestamp 1644511149
transform 1 0 22540 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_245
timestamp 1644511149
transform 1 0 23644 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_251
timestamp 1644511149
transform 1 0 24196 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_90_253
timestamp 1644511149
transform 1 0 24380 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_265
timestamp 1644511149
transform 1 0 25484 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_277
timestamp 1644511149
transform 1 0 26588 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_289
timestamp 1644511149
transform 1 0 27692 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_301
timestamp 1644511149
transform 1 0 28796 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_307
timestamp 1644511149
transform 1 0 29348 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_90_309
timestamp 1644511149
transform 1 0 29532 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_321
timestamp 1644511149
transform 1 0 30636 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_333
timestamp 1644511149
transform 1 0 31740 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_345
timestamp 1644511149
transform 1 0 32844 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_357
timestamp 1644511149
transform 1 0 33948 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_363
timestamp 1644511149
transform 1 0 34500 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_90_365
timestamp 1644511149
transform 1 0 34684 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_377
timestamp 1644511149
transform 1 0 35788 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_389
timestamp 1644511149
transform 1 0 36892 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_401
timestamp 1644511149
transform 1 0 37996 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_413
timestamp 1644511149
transform 1 0 39100 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_419
timestamp 1644511149
transform 1 0 39652 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_90_421
timestamp 1644511149
transform 1 0 39836 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_433
timestamp 1644511149
transform 1 0 40940 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_445
timestamp 1644511149
transform 1 0 42044 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_457
timestamp 1644511149
transform 1 0 43148 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_469
timestamp 1644511149
transform 1 0 44252 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_475
timestamp 1644511149
transform 1 0 44804 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_90_477
timestamp 1644511149
transform 1 0 44988 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_489
timestamp 1644511149
transform 1 0 46092 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_501
timestamp 1644511149
transform 1 0 47196 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_513
timestamp 1644511149
transform 1 0 48300 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_525
timestamp 1644511149
transform 1 0 49404 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_531
timestamp 1644511149
transform 1 0 49956 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_90_533
timestamp 1644511149
transform 1 0 50140 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_545
timestamp 1644511149
transform 1 0 51244 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_557
timestamp 1644511149
transform 1 0 52348 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_569
timestamp 1644511149
transform 1 0 53452 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_581
timestamp 1644511149
transform 1 0 54556 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_587
timestamp 1644511149
transform 1 0 55108 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_90_589
timestamp 1644511149
transform 1 0 55292 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_601
timestamp 1644511149
transform 1 0 56396 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_613
timestamp 1644511149
transform 1 0 57500 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_625
timestamp 1644511149
transform 1 0 58604 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_637
timestamp 1644511149
transform 1 0 59708 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_643
timestamp 1644511149
transform 1 0 60260 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_90_645
timestamp 1644511149
transform 1 0 60444 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_657
timestamp 1644511149
transform 1 0 61548 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_669
timestamp 1644511149
transform 1 0 62652 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_681
timestamp 1644511149
transform 1 0 63756 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_693
timestamp 1644511149
transform 1 0 64860 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_699
timestamp 1644511149
transform 1 0 65412 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_90_701
timestamp 1644511149
transform 1 0 65596 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_713
timestamp 1644511149
transform 1 0 66700 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_725
timestamp 1644511149
transform 1 0 67804 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_737
timestamp 1644511149
transform 1 0 68908 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_749
timestamp 1644511149
transform 1 0 70012 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_755
timestamp 1644511149
transform 1 0 70564 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_90_757
timestamp 1644511149
transform 1 0 70748 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_769
timestamp 1644511149
transform 1 0 71852 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_781
timestamp 1644511149
transform 1 0 72956 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_793
timestamp 1644511149
transform 1 0 74060 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_805
timestamp 1644511149
transform 1 0 75164 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_811
timestamp 1644511149
transform 1 0 75716 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_90_813
timestamp 1644511149
transform 1 0 75900 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_825
timestamp 1644511149
transform 1 0 77004 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_90_837
timestamp 1644511149
transform 1 0 78108 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_90_841
timestamp 1644511149
transform 1 0 78476 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_91_3
timestamp 1644511149
transform 1 0 1380 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_15
timestamp 1644511149
transform 1 0 2484 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_27
timestamp 1644511149
transform 1 0 3588 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_39
timestamp 1644511149
transform 1 0 4692 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_91_51
timestamp 1644511149
transform 1 0 5796 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_91_55
timestamp 1644511149
transform 1 0 6164 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_91_57
timestamp 1644511149
transform 1 0 6348 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_69
timestamp 1644511149
transform 1 0 7452 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_81
timestamp 1644511149
transform 1 0 8556 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_93
timestamp 1644511149
transform 1 0 9660 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_105
timestamp 1644511149
transform 1 0 10764 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_111
timestamp 1644511149
transform 1 0 11316 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_91_113
timestamp 1644511149
transform 1 0 11500 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_125
timestamp 1644511149
transform 1 0 12604 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_137
timestamp 1644511149
transform 1 0 13708 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_149
timestamp 1644511149
transform 1 0 14812 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_161
timestamp 1644511149
transform 1 0 15916 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_167
timestamp 1644511149
transform 1 0 16468 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_91_169
timestamp 1644511149
transform 1 0 16652 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_181
timestamp 1644511149
transform 1 0 17756 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_193
timestamp 1644511149
transform 1 0 18860 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_205
timestamp 1644511149
transform 1 0 19964 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_217
timestamp 1644511149
transform 1 0 21068 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_223
timestamp 1644511149
transform 1 0 21620 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_91_225
timestamp 1644511149
transform 1 0 21804 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_237
timestamp 1644511149
transform 1 0 22908 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_249
timestamp 1644511149
transform 1 0 24012 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_261
timestamp 1644511149
transform 1 0 25116 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_273
timestamp 1644511149
transform 1 0 26220 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_279
timestamp 1644511149
transform 1 0 26772 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_91_281
timestamp 1644511149
transform 1 0 26956 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_293
timestamp 1644511149
transform 1 0 28060 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_305
timestamp 1644511149
transform 1 0 29164 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_317
timestamp 1644511149
transform 1 0 30268 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_329
timestamp 1644511149
transform 1 0 31372 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_335
timestamp 1644511149
transform 1 0 31924 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_91_337
timestamp 1644511149
transform 1 0 32108 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_349
timestamp 1644511149
transform 1 0 33212 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_361
timestamp 1644511149
transform 1 0 34316 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_373
timestamp 1644511149
transform 1 0 35420 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_385
timestamp 1644511149
transform 1 0 36524 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_391
timestamp 1644511149
transform 1 0 37076 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_91_393
timestamp 1644511149
transform 1 0 37260 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_405
timestamp 1644511149
transform 1 0 38364 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_417
timestamp 1644511149
transform 1 0 39468 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_429
timestamp 1644511149
transform 1 0 40572 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_441
timestamp 1644511149
transform 1 0 41676 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_447
timestamp 1644511149
transform 1 0 42228 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_91_449
timestamp 1644511149
transform 1 0 42412 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_461
timestamp 1644511149
transform 1 0 43516 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_473
timestamp 1644511149
transform 1 0 44620 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_485
timestamp 1644511149
transform 1 0 45724 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_497
timestamp 1644511149
transform 1 0 46828 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_503
timestamp 1644511149
transform 1 0 47380 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_91_505
timestamp 1644511149
transform 1 0 47564 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_517
timestamp 1644511149
transform 1 0 48668 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_529
timestamp 1644511149
transform 1 0 49772 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_541
timestamp 1644511149
transform 1 0 50876 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_553
timestamp 1644511149
transform 1 0 51980 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_559
timestamp 1644511149
transform 1 0 52532 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_91_561
timestamp 1644511149
transform 1 0 52716 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_573
timestamp 1644511149
transform 1 0 53820 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_585
timestamp 1644511149
transform 1 0 54924 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_597
timestamp 1644511149
transform 1 0 56028 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_609
timestamp 1644511149
transform 1 0 57132 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_615
timestamp 1644511149
transform 1 0 57684 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_91_617
timestamp 1644511149
transform 1 0 57868 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_629
timestamp 1644511149
transform 1 0 58972 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_641
timestamp 1644511149
transform 1 0 60076 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_653
timestamp 1644511149
transform 1 0 61180 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_665
timestamp 1644511149
transform 1 0 62284 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_671
timestamp 1644511149
transform 1 0 62836 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_91_673
timestamp 1644511149
transform 1 0 63020 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_685
timestamp 1644511149
transform 1 0 64124 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_697
timestamp 1644511149
transform 1 0 65228 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_709
timestamp 1644511149
transform 1 0 66332 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_721
timestamp 1644511149
transform 1 0 67436 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_727
timestamp 1644511149
transform 1 0 67988 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_91_729
timestamp 1644511149
transform 1 0 68172 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_741
timestamp 1644511149
transform 1 0 69276 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_753
timestamp 1644511149
transform 1 0 70380 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_765
timestamp 1644511149
transform 1 0 71484 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_777
timestamp 1644511149
transform 1 0 72588 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_783
timestamp 1644511149
transform 1 0 73140 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_91_785
timestamp 1644511149
transform 1 0 73324 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_797
timestamp 1644511149
transform 1 0 74428 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_809
timestamp 1644511149
transform 1 0 75532 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_91_821
timestamp 1644511149
transform 1 0 76636 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_91_829
timestamp 1644511149
transform 1 0 77372 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_91_836
timestamp 1644511149
transform 1 0 78016 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_91_841
timestamp 1644511149
transform 1 0 78476 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_92_3
timestamp 1644511149
transform 1 0 1380 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_15
timestamp 1644511149
transform 1 0 2484 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_92_27
timestamp 1644511149
transform 1 0 3588 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_92_29
timestamp 1644511149
transform 1 0 3772 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_41
timestamp 1644511149
transform 1 0 4876 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_53
timestamp 1644511149
transform 1 0 5980 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_65
timestamp 1644511149
transform 1 0 7084 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_77
timestamp 1644511149
transform 1 0 8188 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_83
timestamp 1644511149
transform 1 0 8740 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_92_85
timestamp 1644511149
transform 1 0 8924 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_97
timestamp 1644511149
transform 1 0 10028 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_109
timestamp 1644511149
transform 1 0 11132 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_121
timestamp 1644511149
transform 1 0 12236 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_133
timestamp 1644511149
transform 1 0 13340 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_139
timestamp 1644511149
transform 1 0 13892 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_92_141
timestamp 1644511149
transform 1 0 14076 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_153
timestamp 1644511149
transform 1 0 15180 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_165
timestamp 1644511149
transform 1 0 16284 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_177
timestamp 1644511149
transform 1 0 17388 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_189
timestamp 1644511149
transform 1 0 18492 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_195
timestamp 1644511149
transform 1 0 19044 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_92_197
timestamp 1644511149
transform 1 0 19228 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_209
timestamp 1644511149
transform 1 0 20332 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_221
timestamp 1644511149
transform 1 0 21436 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_233
timestamp 1644511149
transform 1 0 22540 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_245
timestamp 1644511149
transform 1 0 23644 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_251
timestamp 1644511149
transform 1 0 24196 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_92_253
timestamp 1644511149
transform 1 0 24380 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_265
timestamp 1644511149
transform 1 0 25484 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_277
timestamp 1644511149
transform 1 0 26588 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_289
timestamp 1644511149
transform 1 0 27692 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_301
timestamp 1644511149
transform 1 0 28796 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_307
timestamp 1644511149
transform 1 0 29348 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_92_309
timestamp 1644511149
transform 1 0 29532 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_321
timestamp 1644511149
transform 1 0 30636 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_333
timestamp 1644511149
transform 1 0 31740 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_345
timestamp 1644511149
transform 1 0 32844 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_357
timestamp 1644511149
transform 1 0 33948 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_363
timestamp 1644511149
transform 1 0 34500 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_92_365
timestamp 1644511149
transform 1 0 34684 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_377
timestamp 1644511149
transform 1 0 35788 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_389
timestamp 1644511149
transform 1 0 36892 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_401
timestamp 1644511149
transform 1 0 37996 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_413
timestamp 1644511149
transform 1 0 39100 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_419
timestamp 1644511149
transform 1 0 39652 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_92_421
timestamp 1644511149
transform 1 0 39836 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_433
timestamp 1644511149
transform 1 0 40940 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_445
timestamp 1644511149
transform 1 0 42044 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_457
timestamp 1644511149
transform 1 0 43148 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_469
timestamp 1644511149
transform 1 0 44252 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_475
timestamp 1644511149
transform 1 0 44804 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_92_477
timestamp 1644511149
transform 1 0 44988 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_489
timestamp 1644511149
transform 1 0 46092 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_501
timestamp 1644511149
transform 1 0 47196 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_513
timestamp 1644511149
transform 1 0 48300 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_525
timestamp 1644511149
transform 1 0 49404 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_531
timestamp 1644511149
transform 1 0 49956 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_92_533
timestamp 1644511149
transform 1 0 50140 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_545
timestamp 1644511149
transform 1 0 51244 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_557
timestamp 1644511149
transform 1 0 52348 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_569
timestamp 1644511149
transform 1 0 53452 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_581
timestamp 1644511149
transform 1 0 54556 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_587
timestamp 1644511149
transform 1 0 55108 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_92_589
timestamp 1644511149
transform 1 0 55292 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_601
timestamp 1644511149
transform 1 0 56396 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_613
timestamp 1644511149
transform 1 0 57500 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_625
timestamp 1644511149
transform 1 0 58604 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_637
timestamp 1644511149
transform 1 0 59708 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_643
timestamp 1644511149
transform 1 0 60260 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_92_645
timestamp 1644511149
transform 1 0 60444 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_657
timestamp 1644511149
transform 1 0 61548 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_669
timestamp 1644511149
transform 1 0 62652 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_681
timestamp 1644511149
transform 1 0 63756 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_693
timestamp 1644511149
transform 1 0 64860 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_699
timestamp 1644511149
transform 1 0 65412 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_92_701
timestamp 1644511149
transform 1 0 65596 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_713
timestamp 1644511149
transform 1 0 66700 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_725
timestamp 1644511149
transform 1 0 67804 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_737
timestamp 1644511149
transform 1 0 68908 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_749
timestamp 1644511149
transform 1 0 70012 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_755
timestamp 1644511149
transform 1 0 70564 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_92_757
timestamp 1644511149
transform 1 0 70748 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_769
timestamp 1644511149
transform 1 0 71852 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_781
timestamp 1644511149
transform 1 0 72956 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_793
timestamp 1644511149
transform 1 0 74060 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_805
timestamp 1644511149
transform 1 0 75164 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_811
timestamp 1644511149
transform 1 0 75716 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_92_813
timestamp 1644511149
transform 1 0 75900 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_825
timestamp 1644511149
transform 1 0 77004 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_92_837
timestamp 1644511149
transform 1 0 78108 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_92_841
timestamp 1644511149
transform 1 0 78476 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_93_3
timestamp 1644511149
transform 1 0 1380 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_15
timestamp 1644511149
transform 1 0 2484 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_27
timestamp 1644511149
transform 1 0 3588 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_39
timestamp 1644511149
transform 1 0 4692 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_93_51
timestamp 1644511149
transform 1 0 5796 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_93_55
timestamp 1644511149
transform 1 0 6164 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_93_57
timestamp 1644511149
transform 1 0 6348 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_69
timestamp 1644511149
transform 1 0 7452 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_81
timestamp 1644511149
transform 1 0 8556 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_93
timestamp 1644511149
transform 1 0 9660 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_105
timestamp 1644511149
transform 1 0 10764 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_111
timestamp 1644511149
transform 1 0 11316 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_93_113
timestamp 1644511149
transform 1 0 11500 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_125
timestamp 1644511149
transform 1 0 12604 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_137
timestamp 1644511149
transform 1 0 13708 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_149
timestamp 1644511149
transform 1 0 14812 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_161
timestamp 1644511149
transform 1 0 15916 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_167
timestamp 1644511149
transform 1 0 16468 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_93_169
timestamp 1644511149
transform 1 0 16652 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_181
timestamp 1644511149
transform 1 0 17756 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_193
timestamp 1644511149
transform 1 0 18860 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_205
timestamp 1644511149
transform 1 0 19964 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_217
timestamp 1644511149
transform 1 0 21068 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_223
timestamp 1644511149
transform 1 0 21620 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_93_225
timestamp 1644511149
transform 1 0 21804 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_237
timestamp 1644511149
transform 1 0 22908 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_249
timestamp 1644511149
transform 1 0 24012 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_261
timestamp 1644511149
transform 1 0 25116 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_273
timestamp 1644511149
transform 1 0 26220 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_279
timestamp 1644511149
transform 1 0 26772 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_93_281
timestamp 1644511149
transform 1 0 26956 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_293
timestamp 1644511149
transform 1 0 28060 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_305
timestamp 1644511149
transform 1 0 29164 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_317
timestamp 1644511149
transform 1 0 30268 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_329
timestamp 1644511149
transform 1 0 31372 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_335
timestamp 1644511149
transform 1 0 31924 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_93_337
timestamp 1644511149
transform 1 0 32108 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_349
timestamp 1644511149
transform 1 0 33212 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_361
timestamp 1644511149
transform 1 0 34316 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_373
timestamp 1644511149
transform 1 0 35420 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_385
timestamp 1644511149
transform 1 0 36524 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_391
timestamp 1644511149
transform 1 0 37076 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_93_393
timestamp 1644511149
transform 1 0 37260 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_405
timestamp 1644511149
transform 1 0 38364 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_417
timestamp 1644511149
transform 1 0 39468 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_429
timestamp 1644511149
transform 1 0 40572 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_441
timestamp 1644511149
transform 1 0 41676 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_447
timestamp 1644511149
transform 1 0 42228 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_93_449
timestamp 1644511149
transform 1 0 42412 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_461
timestamp 1644511149
transform 1 0 43516 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_473
timestamp 1644511149
transform 1 0 44620 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_485
timestamp 1644511149
transform 1 0 45724 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_497
timestamp 1644511149
transform 1 0 46828 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_503
timestamp 1644511149
transform 1 0 47380 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_93_505
timestamp 1644511149
transform 1 0 47564 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_517
timestamp 1644511149
transform 1 0 48668 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_529
timestamp 1644511149
transform 1 0 49772 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_541
timestamp 1644511149
transform 1 0 50876 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_553
timestamp 1644511149
transform 1 0 51980 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_559
timestamp 1644511149
transform 1 0 52532 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_93_561
timestamp 1644511149
transform 1 0 52716 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_573
timestamp 1644511149
transform 1 0 53820 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_585
timestamp 1644511149
transform 1 0 54924 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_597
timestamp 1644511149
transform 1 0 56028 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_609
timestamp 1644511149
transform 1 0 57132 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_615
timestamp 1644511149
transform 1 0 57684 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_93_617
timestamp 1644511149
transform 1 0 57868 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_629
timestamp 1644511149
transform 1 0 58972 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_641
timestamp 1644511149
transform 1 0 60076 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_653
timestamp 1644511149
transform 1 0 61180 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_665
timestamp 1644511149
transform 1 0 62284 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_671
timestamp 1644511149
transform 1 0 62836 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_93_673
timestamp 1644511149
transform 1 0 63020 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_685
timestamp 1644511149
transform 1 0 64124 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_697
timestamp 1644511149
transform 1 0 65228 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_709
timestamp 1644511149
transform 1 0 66332 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_721
timestamp 1644511149
transform 1 0 67436 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_727
timestamp 1644511149
transform 1 0 67988 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_93_729
timestamp 1644511149
transform 1 0 68172 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_741
timestamp 1644511149
transform 1 0 69276 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_753
timestamp 1644511149
transform 1 0 70380 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_765
timestamp 1644511149
transform 1 0 71484 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_777
timestamp 1644511149
transform 1 0 72588 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_783
timestamp 1644511149
transform 1 0 73140 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_93_785
timestamp 1644511149
transform 1 0 73324 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_797
timestamp 1644511149
transform 1 0 74428 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_809
timestamp 1644511149
transform 1 0 75532 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_821
timestamp 1644511149
transform 1 0 76636 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_833
timestamp 1644511149
transform 1 0 77740 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_839
timestamp 1644511149
transform 1 0 78292 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_93_841
timestamp 1644511149
transform 1 0 78476 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_94_3
timestamp 1644511149
transform 1 0 1380 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_15
timestamp 1644511149
transform 1 0 2484 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_94_27
timestamp 1644511149
transform 1 0 3588 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_94_29
timestamp 1644511149
transform 1 0 3772 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_41
timestamp 1644511149
transform 1 0 4876 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_53
timestamp 1644511149
transform 1 0 5980 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_65
timestamp 1644511149
transform 1 0 7084 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_77
timestamp 1644511149
transform 1 0 8188 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_83
timestamp 1644511149
transform 1 0 8740 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_94_85
timestamp 1644511149
transform 1 0 8924 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_97
timestamp 1644511149
transform 1 0 10028 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_109
timestamp 1644511149
transform 1 0 11132 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_121
timestamp 1644511149
transform 1 0 12236 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_133
timestamp 1644511149
transform 1 0 13340 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_139
timestamp 1644511149
transform 1 0 13892 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_94_141
timestamp 1644511149
transform 1 0 14076 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_153
timestamp 1644511149
transform 1 0 15180 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_165
timestamp 1644511149
transform 1 0 16284 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_177
timestamp 1644511149
transform 1 0 17388 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_189
timestamp 1644511149
transform 1 0 18492 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_195
timestamp 1644511149
transform 1 0 19044 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_94_197
timestamp 1644511149
transform 1 0 19228 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_209
timestamp 1644511149
transform 1 0 20332 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_221
timestamp 1644511149
transform 1 0 21436 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_233
timestamp 1644511149
transform 1 0 22540 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_245
timestamp 1644511149
transform 1 0 23644 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_251
timestamp 1644511149
transform 1 0 24196 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_94_253
timestamp 1644511149
transform 1 0 24380 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_265
timestamp 1644511149
transform 1 0 25484 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_277
timestamp 1644511149
transform 1 0 26588 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_289
timestamp 1644511149
transform 1 0 27692 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_301
timestamp 1644511149
transform 1 0 28796 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_307
timestamp 1644511149
transform 1 0 29348 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_94_309
timestamp 1644511149
transform 1 0 29532 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_321
timestamp 1644511149
transform 1 0 30636 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_333
timestamp 1644511149
transform 1 0 31740 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_345
timestamp 1644511149
transform 1 0 32844 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_357
timestamp 1644511149
transform 1 0 33948 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_363
timestamp 1644511149
transform 1 0 34500 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_94_365
timestamp 1644511149
transform 1 0 34684 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_377
timestamp 1644511149
transform 1 0 35788 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_389
timestamp 1644511149
transform 1 0 36892 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_401
timestamp 1644511149
transform 1 0 37996 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_413
timestamp 1644511149
transform 1 0 39100 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_419
timestamp 1644511149
transform 1 0 39652 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_94_421
timestamp 1644511149
transform 1 0 39836 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_433
timestamp 1644511149
transform 1 0 40940 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_445
timestamp 1644511149
transform 1 0 42044 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_457
timestamp 1644511149
transform 1 0 43148 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_469
timestamp 1644511149
transform 1 0 44252 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_475
timestamp 1644511149
transform 1 0 44804 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_94_477
timestamp 1644511149
transform 1 0 44988 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_489
timestamp 1644511149
transform 1 0 46092 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_501
timestamp 1644511149
transform 1 0 47196 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_513
timestamp 1644511149
transform 1 0 48300 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_525
timestamp 1644511149
transform 1 0 49404 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_531
timestamp 1644511149
transform 1 0 49956 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_94_533
timestamp 1644511149
transform 1 0 50140 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_545
timestamp 1644511149
transform 1 0 51244 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_557
timestamp 1644511149
transform 1 0 52348 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_569
timestamp 1644511149
transform 1 0 53452 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_581
timestamp 1644511149
transform 1 0 54556 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_587
timestamp 1644511149
transform 1 0 55108 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_94_589
timestamp 1644511149
transform 1 0 55292 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_601
timestamp 1644511149
transform 1 0 56396 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_613
timestamp 1644511149
transform 1 0 57500 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_625
timestamp 1644511149
transform 1 0 58604 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_637
timestamp 1644511149
transform 1 0 59708 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_643
timestamp 1644511149
transform 1 0 60260 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_94_645
timestamp 1644511149
transform 1 0 60444 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_657
timestamp 1644511149
transform 1 0 61548 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_669
timestamp 1644511149
transform 1 0 62652 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_681
timestamp 1644511149
transform 1 0 63756 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_693
timestamp 1644511149
transform 1 0 64860 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_699
timestamp 1644511149
transform 1 0 65412 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_94_701
timestamp 1644511149
transform 1 0 65596 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_713
timestamp 1644511149
transform 1 0 66700 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_725
timestamp 1644511149
transform 1 0 67804 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_737
timestamp 1644511149
transform 1 0 68908 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_749
timestamp 1644511149
transform 1 0 70012 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_755
timestamp 1644511149
transform 1 0 70564 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_94_757
timestamp 1644511149
transform 1 0 70748 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_769
timestamp 1644511149
transform 1 0 71852 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_781
timestamp 1644511149
transform 1 0 72956 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_793
timestamp 1644511149
transform 1 0 74060 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_805
timestamp 1644511149
transform 1 0 75164 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_811
timestamp 1644511149
transform 1 0 75716 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_94_813
timestamp 1644511149
transform 1 0 75900 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_825
timestamp 1644511149
transform 1 0 77004 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_94_837
timestamp 1644511149
transform 1 0 78108 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_94_841
timestamp 1644511149
transform 1 0 78476 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_95_3
timestamp 1644511149
transform 1 0 1380 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_15
timestamp 1644511149
transform 1 0 2484 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_27
timestamp 1644511149
transform 1 0 3588 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_39
timestamp 1644511149
transform 1 0 4692 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_95_51
timestamp 1644511149
transform 1 0 5796 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_95_55
timestamp 1644511149
transform 1 0 6164 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_95_57
timestamp 1644511149
transform 1 0 6348 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_69
timestamp 1644511149
transform 1 0 7452 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_81
timestamp 1644511149
transform 1 0 8556 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_93
timestamp 1644511149
transform 1 0 9660 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_105
timestamp 1644511149
transform 1 0 10764 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_111
timestamp 1644511149
transform 1 0 11316 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_95_113
timestamp 1644511149
transform 1 0 11500 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_125
timestamp 1644511149
transform 1 0 12604 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_137
timestamp 1644511149
transform 1 0 13708 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_149
timestamp 1644511149
transform 1 0 14812 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_161
timestamp 1644511149
transform 1 0 15916 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_167
timestamp 1644511149
transform 1 0 16468 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_95_169
timestamp 1644511149
transform 1 0 16652 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_181
timestamp 1644511149
transform 1 0 17756 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_193
timestamp 1644511149
transform 1 0 18860 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_205
timestamp 1644511149
transform 1 0 19964 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_217
timestamp 1644511149
transform 1 0 21068 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_223
timestamp 1644511149
transform 1 0 21620 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_95_225
timestamp 1644511149
transform 1 0 21804 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_237
timestamp 1644511149
transform 1 0 22908 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_249
timestamp 1644511149
transform 1 0 24012 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_261
timestamp 1644511149
transform 1 0 25116 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_273
timestamp 1644511149
transform 1 0 26220 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_279
timestamp 1644511149
transform 1 0 26772 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_95_281
timestamp 1644511149
transform 1 0 26956 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_293
timestamp 1644511149
transform 1 0 28060 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_305
timestamp 1644511149
transform 1 0 29164 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_317
timestamp 1644511149
transform 1 0 30268 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_329
timestamp 1644511149
transform 1 0 31372 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_335
timestamp 1644511149
transform 1 0 31924 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_95_337
timestamp 1644511149
transform 1 0 32108 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_349
timestamp 1644511149
transform 1 0 33212 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_361
timestamp 1644511149
transform 1 0 34316 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_373
timestamp 1644511149
transform 1 0 35420 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_385
timestamp 1644511149
transform 1 0 36524 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_391
timestamp 1644511149
transform 1 0 37076 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_95_393
timestamp 1644511149
transform 1 0 37260 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_405
timestamp 1644511149
transform 1 0 38364 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_417
timestamp 1644511149
transform 1 0 39468 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_429
timestamp 1644511149
transform 1 0 40572 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_441
timestamp 1644511149
transform 1 0 41676 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_447
timestamp 1644511149
transform 1 0 42228 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_95_449
timestamp 1644511149
transform 1 0 42412 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_461
timestamp 1644511149
transform 1 0 43516 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_473
timestamp 1644511149
transform 1 0 44620 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_485
timestamp 1644511149
transform 1 0 45724 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_497
timestamp 1644511149
transform 1 0 46828 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_503
timestamp 1644511149
transform 1 0 47380 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_95_505
timestamp 1644511149
transform 1 0 47564 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_517
timestamp 1644511149
transform 1 0 48668 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_529
timestamp 1644511149
transform 1 0 49772 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_541
timestamp 1644511149
transform 1 0 50876 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_553
timestamp 1644511149
transform 1 0 51980 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_559
timestamp 1644511149
transform 1 0 52532 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_95_561
timestamp 1644511149
transform 1 0 52716 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_573
timestamp 1644511149
transform 1 0 53820 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_585
timestamp 1644511149
transform 1 0 54924 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_597
timestamp 1644511149
transform 1 0 56028 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_609
timestamp 1644511149
transform 1 0 57132 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_615
timestamp 1644511149
transform 1 0 57684 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_95_617
timestamp 1644511149
transform 1 0 57868 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_629
timestamp 1644511149
transform 1 0 58972 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_641
timestamp 1644511149
transform 1 0 60076 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_653
timestamp 1644511149
transform 1 0 61180 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_665
timestamp 1644511149
transform 1 0 62284 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_671
timestamp 1644511149
transform 1 0 62836 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_95_673
timestamp 1644511149
transform 1 0 63020 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_685
timestamp 1644511149
transform 1 0 64124 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_697
timestamp 1644511149
transform 1 0 65228 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_709
timestamp 1644511149
transform 1 0 66332 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_721
timestamp 1644511149
transform 1 0 67436 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_727
timestamp 1644511149
transform 1 0 67988 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_95_729
timestamp 1644511149
transform 1 0 68172 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_741
timestamp 1644511149
transform 1 0 69276 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_753
timestamp 1644511149
transform 1 0 70380 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_765
timestamp 1644511149
transform 1 0 71484 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_777
timestamp 1644511149
transform 1 0 72588 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_783
timestamp 1644511149
transform 1 0 73140 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_95_785
timestamp 1644511149
transform 1 0 73324 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_797
timestamp 1644511149
transform 1 0 74428 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_809
timestamp 1644511149
transform 1 0 75532 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_821
timestamp 1644511149
transform 1 0 76636 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_833
timestamp 1644511149
transform 1 0 77740 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_839
timestamp 1644511149
transform 1 0 78292 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_95_841
timestamp 1644511149
transform 1 0 78476 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_96_7
timestamp 1644511149
transform 1 0 1748 0 1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_96_11
timestamp 1644511149
transform 1 0 2116 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_96_23
timestamp 1644511149
transform 1 0 3220 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_96_27
timestamp 1644511149
transform 1 0 3588 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_96_29
timestamp 1644511149
transform 1 0 3772 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_41
timestamp 1644511149
transform 1 0 4876 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_53
timestamp 1644511149
transform 1 0 5980 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_65
timestamp 1644511149
transform 1 0 7084 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_77
timestamp 1644511149
transform 1 0 8188 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_83
timestamp 1644511149
transform 1 0 8740 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_96_85
timestamp 1644511149
transform 1 0 8924 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_97
timestamp 1644511149
transform 1 0 10028 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_109
timestamp 1644511149
transform 1 0 11132 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_121
timestamp 1644511149
transform 1 0 12236 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_133
timestamp 1644511149
transform 1 0 13340 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_139
timestamp 1644511149
transform 1 0 13892 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_96_141
timestamp 1644511149
transform 1 0 14076 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_153
timestamp 1644511149
transform 1 0 15180 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_165
timestamp 1644511149
transform 1 0 16284 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_177
timestamp 1644511149
transform 1 0 17388 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_189
timestamp 1644511149
transform 1 0 18492 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_195
timestamp 1644511149
transform 1 0 19044 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_96_197
timestamp 1644511149
transform 1 0 19228 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_209
timestamp 1644511149
transform 1 0 20332 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_221
timestamp 1644511149
transform 1 0 21436 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_233
timestamp 1644511149
transform 1 0 22540 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_245
timestamp 1644511149
transform 1 0 23644 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_251
timestamp 1644511149
transform 1 0 24196 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_96_253
timestamp 1644511149
transform 1 0 24380 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_265
timestamp 1644511149
transform 1 0 25484 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_277
timestamp 1644511149
transform 1 0 26588 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_289
timestamp 1644511149
transform 1 0 27692 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_301
timestamp 1644511149
transform 1 0 28796 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_307
timestamp 1644511149
transform 1 0 29348 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_96_309
timestamp 1644511149
transform 1 0 29532 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_321
timestamp 1644511149
transform 1 0 30636 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_333
timestamp 1644511149
transform 1 0 31740 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_345
timestamp 1644511149
transform 1 0 32844 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_357
timestamp 1644511149
transform 1 0 33948 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_363
timestamp 1644511149
transform 1 0 34500 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_96_365
timestamp 1644511149
transform 1 0 34684 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_377
timestamp 1644511149
transform 1 0 35788 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_389
timestamp 1644511149
transform 1 0 36892 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_401
timestamp 1644511149
transform 1 0 37996 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_413
timestamp 1644511149
transform 1 0 39100 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_419
timestamp 1644511149
transform 1 0 39652 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_96_421
timestamp 1644511149
transform 1 0 39836 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_433
timestamp 1644511149
transform 1 0 40940 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_445
timestamp 1644511149
transform 1 0 42044 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_457
timestamp 1644511149
transform 1 0 43148 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_469
timestamp 1644511149
transform 1 0 44252 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_475
timestamp 1644511149
transform 1 0 44804 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_96_477
timestamp 1644511149
transform 1 0 44988 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_489
timestamp 1644511149
transform 1 0 46092 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_501
timestamp 1644511149
transform 1 0 47196 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_513
timestamp 1644511149
transform 1 0 48300 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_525
timestamp 1644511149
transform 1 0 49404 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_531
timestamp 1644511149
transform 1 0 49956 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_96_533
timestamp 1644511149
transform 1 0 50140 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_545
timestamp 1644511149
transform 1 0 51244 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_557
timestamp 1644511149
transform 1 0 52348 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_569
timestamp 1644511149
transform 1 0 53452 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_581
timestamp 1644511149
transform 1 0 54556 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_587
timestamp 1644511149
transform 1 0 55108 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_96_589
timestamp 1644511149
transform 1 0 55292 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_601
timestamp 1644511149
transform 1 0 56396 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_613
timestamp 1644511149
transform 1 0 57500 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_625
timestamp 1644511149
transform 1 0 58604 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_637
timestamp 1644511149
transform 1 0 59708 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_643
timestamp 1644511149
transform 1 0 60260 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_96_645
timestamp 1644511149
transform 1 0 60444 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_657
timestamp 1644511149
transform 1 0 61548 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_669
timestamp 1644511149
transform 1 0 62652 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_681
timestamp 1644511149
transform 1 0 63756 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_693
timestamp 1644511149
transform 1 0 64860 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_699
timestamp 1644511149
transform 1 0 65412 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_96_701
timestamp 1644511149
transform 1 0 65596 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_713
timestamp 1644511149
transform 1 0 66700 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_725
timestamp 1644511149
transform 1 0 67804 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_737
timestamp 1644511149
transform 1 0 68908 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_749
timestamp 1644511149
transform 1 0 70012 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_755
timestamp 1644511149
transform 1 0 70564 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_96_757
timestamp 1644511149
transform 1 0 70748 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_769
timestamp 1644511149
transform 1 0 71852 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_781
timestamp 1644511149
transform 1 0 72956 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_793
timestamp 1644511149
transform 1 0 74060 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_805
timestamp 1644511149
transform 1 0 75164 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_811
timestamp 1644511149
transform 1 0 75716 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_96_813
timestamp 1644511149
transform 1 0 75900 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_825
timestamp 1644511149
transform 1 0 77004 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_96_837
timestamp 1644511149
transform 1 0 78108 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_96_841
timestamp 1644511149
transform 1 0 78476 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_97_3
timestamp 1644511149
transform 1 0 1380 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_15
timestamp 1644511149
transform 1 0 2484 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_27
timestamp 1644511149
transform 1 0 3588 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_39
timestamp 1644511149
transform 1 0 4692 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_97_51
timestamp 1644511149
transform 1 0 5796 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_97_55
timestamp 1644511149
transform 1 0 6164 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_97_57
timestamp 1644511149
transform 1 0 6348 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_69
timestamp 1644511149
transform 1 0 7452 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_81
timestamp 1644511149
transform 1 0 8556 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_93
timestamp 1644511149
transform 1 0 9660 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_105
timestamp 1644511149
transform 1 0 10764 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_111
timestamp 1644511149
transform 1 0 11316 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_97_113
timestamp 1644511149
transform 1 0 11500 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_125
timestamp 1644511149
transform 1 0 12604 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_137
timestamp 1644511149
transform 1 0 13708 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_149
timestamp 1644511149
transform 1 0 14812 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_161
timestamp 1644511149
transform 1 0 15916 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_167
timestamp 1644511149
transform 1 0 16468 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_97_169
timestamp 1644511149
transform 1 0 16652 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_181
timestamp 1644511149
transform 1 0 17756 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_193
timestamp 1644511149
transform 1 0 18860 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_205
timestamp 1644511149
transform 1 0 19964 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_217
timestamp 1644511149
transform 1 0 21068 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_223
timestamp 1644511149
transform 1 0 21620 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_97_225
timestamp 1644511149
transform 1 0 21804 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_237
timestamp 1644511149
transform 1 0 22908 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_249
timestamp 1644511149
transform 1 0 24012 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_261
timestamp 1644511149
transform 1 0 25116 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_273
timestamp 1644511149
transform 1 0 26220 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_279
timestamp 1644511149
transform 1 0 26772 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_97_281
timestamp 1644511149
transform 1 0 26956 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_293
timestamp 1644511149
transform 1 0 28060 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_305
timestamp 1644511149
transform 1 0 29164 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_317
timestamp 1644511149
transform 1 0 30268 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_329
timestamp 1644511149
transform 1 0 31372 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_335
timestamp 1644511149
transform 1 0 31924 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_97_337
timestamp 1644511149
transform 1 0 32108 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_349
timestamp 1644511149
transform 1 0 33212 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_361
timestamp 1644511149
transform 1 0 34316 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_373
timestamp 1644511149
transform 1 0 35420 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_385
timestamp 1644511149
transform 1 0 36524 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_391
timestamp 1644511149
transform 1 0 37076 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_97_393
timestamp 1644511149
transform 1 0 37260 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_405
timestamp 1644511149
transform 1 0 38364 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_417
timestamp 1644511149
transform 1 0 39468 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_429
timestamp 1644511149
transform 1 0 40572 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_441
timestamp 1644511149
transform 1 0 41676 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_447
timestamp 1644511149
transform 1 0 42228 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_97_449
timestamp 1644511149
transform 1 0 42412 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_461
timestamp 1644511149
transform 1 0 43516 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_473
timestamp 1644511149
transform 1 0 44620 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_485
timestamp 1644511149
transform 1 0 45724 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_497
timestamp 1644511149
transform 1 0 46828 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_503
timestamp 1644511149
transform 1 0 47380 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_97_505
timestamp 1644511149
transform 1 0 47564 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_517
timestamp 1644511149
transform 1 0 48668 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_529
timestamp 1644511149
transform 1 0 49772 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_541
timestamp 1644511149
transform 1 0 50876 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_553
timestamp 1644511149
transform 1 0 51980 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_559
timestamp 1644511149
transform 1 0 52532 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_97_561
timestamp 1644511149
transform 1 0 52716 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_573
timestamp 1644511149
transform 1 0 53820 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_585
timestamp 1644511149
transform 1 0 54924 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_597
timestamp 1644511149
transform 1 0 56028 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_609
timestamp 1644511149
transform 1 0 57132 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_615
timestamp 1644511149
transform 1 0 57684 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_97_617
timestamp 1644511149
transform 1 0 57868 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_629
timestamp 1644511149
transform 1 0 58972 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_641
timestamp 1644511149
transform 1 0 60076 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_653
timestamp 1644511149
transform 1 0 61180 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_665
timestamp 1644511149
transform 1 0 62284 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_671
timestamp 1644511149
transform 1 0 62836 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_97_673
timestamp 1644511149
transform 1 0 63020 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_685
timestamp 1644511149
transform 1 0 64124 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_697
timestamp 1644511149
transform 1 0 65228 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_709
timestamp 1644511149
transform 1 0 66332 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_721
timestamp 1644511149
transform 1 0 67436 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_727
timestamp 1644511149
transform 1 0 67988 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_97_729
timestamp 1644511149
transform 1 0 68172 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_741
timestamp 1644511149
transform 1 0 69276 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_753
timestamp 1644511149
transform 1 0 70380 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_765
timestamp 1644511149
transform 1 0 71484 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_777
timestamp 1644511149
transform 1 0 72588 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_783
timestamp 1644511149
transform 1 0 73140 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_97_785
timestamp 1644511149
transform 1 0 73324 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_797
timestamp 1644511149
transform 1 0 74428 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_809
timestamp 1644511149
transform 1 0 75532 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_821
timestamp 1644511149
transform 1 0 76636 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_833
timestamp 1644511149
transform 1 0 77740 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_839
timestamp 1644511149
transform 1 0 78292 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_97_841
timestamp 1644511149
transform 1 0 78476 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_98_3
timestamp 1644511149
transform 1 0 1380 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_15
timestamp 1644511149
transform 1 0 2484 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_98_27
timestamp 1644511149
transform 1 0 3588 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_98_29
timestamp 1644511149
transform 1 0 3772 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_41
timestamp 1644511149
transform 1 0 4876 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_53
timestamp 1644511149
transform 1 0 5980 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_65
timestamp 1644511149
transform 1 0 7084 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_77
timestamp 1644511149
transform 1 0 8188 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_83
timestamp 1644511149
transform 1 0 8740 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_98_85
timestamp 1644511149
transform 1 0 8924 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_97
timestamp 1644511149
transform 1 0 10028 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_109
timestamp 1644511149
transform 1 0 11132 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_121
timestamp 1644511149
transform 1 0 12236 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_133
timestamp 1644511149
transform 1 0 13340 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_139
timestamp 1644511149
transform 1 0 13892 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_98_141
timestamp 1644511149
transform 1 0 14076 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_153
timestamp 1644511149
transform 1 0 15180 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_165
timestamp 1644511149
transform 1 0 16284 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_177
timestamp 1644511149
transform 1 0 17388 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_189
timestamp 1644511149
transform 1 0 18492 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_195
timestamp 1644511149
transform 1 0 19044 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_98_197
timestamp 1644511149
transform 1 0 19228 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_209
timestamp 1644511149
transform 1 0 20332 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_221
timestamp 1644511149
transform 1 0 21436 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_233
timestamp 1644511149
transform 1 0 22540 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_245
timestamp 1644511149
transform 1 0 23644 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_251
timestamp 1644511149
transform 1 0 24196 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_98_253
timestamp 1644511149
transform 1 0 24380 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_265
timestamp 1644511149
transform 1 0 25484 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_277
timestamp 1644511149
transform 1 0 26588 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_289
timestamp 1644511149
transform 1 0 27692 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_301
timestamp 1644511149
transform 1 0 28796 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_307
timestamp 1644511149
transform 1 0 29348 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_98_309
timestamp 1644511149
transform 1 0 29532 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_321
timestamp 1644511149
transform 1 0 30636 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_333
timestamp 1644511149
transform 1 0 31740 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_345
timestamp 1644511149
transform 1 0 32844 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_357
timestamp 1644511149
transform 1 0 33948 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_363
timestamp 1644511149
transform 1 0 34500 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_98_365
timestamp 1644511149
transform 1 0 34684 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_377
timestamp 1644511149
transform 1 0 35788 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_389
timestamp 1644511149
transform 1 0 36892 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_401
timestamp 1644511149
transform 1 0 37996 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_413
timestamp 1644511149
transform 1 0 39100 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_419
timestamp 1644511149
transform 1 0 39652 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_98_421
timestamp 1644511149
transform 1 0 39836 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_433
timestamp 1644511149
transform 1 0 40940 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_445
timestamp 1644511149
transform 1 0 42044 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_457
timestamp 1644511149
transform 1 0 43148 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_469
timestamp 1644511149
transform 1 0 44252 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_475
timestamp 1644511149
transform 1 0 44804 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_98_477
timestamp 1644511149
transform 1 0 44988 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_489
timestamp 1644511149
transform 1 0 46092 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_501
timestamp 1644511149
transform 1 0 47196 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_513
timestamp 1644511149
transform 1 0 48300 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_525
timestamp 1644511149
transform 1 0 49404 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_531
timestamp 1644511149
transform 1 0 49956 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_98_533
timestamp 1644511149
transform 1 0 50140 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_545
timestamp 1644511149
transform 1 0 51244 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_557
timestamp 1644511149
transform 1 0 52348 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_569
timestamp 1644511149
transform 1 0 53452 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_581
timestamp 1644511149
transform 1 0 54556 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_587
timestamp 1644511149
transform 1 0 55108 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_98_589
timestamp 1644511149
transform 1 0 55292 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_601
timestamp 1644511149
transform 1 0 56396 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_613
timestamp 1644511149
transform 1 0 57500 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_625
timestamp 1644511149
transform 1 0 58604 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_637
timestamp 1644511149
transform 1 0 59708 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_643
timestamp 1644511149
transform 1 0 60260 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_98_645
timestamp 1644511149
transform 1 0 60444 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_657
timestamp 1644511149
transform 1 0 61548 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_669
timestamp 1644511149
transform 1 0 62652 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_681
timestamp 1644511149
transform 1 0 63756 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_693
timestamp 1644511149
transform 1 0 64860 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_699
timestamp 1644511149
transform 1 0 65412 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_98_701
timestamp 1644511149
transform 1 0 65596 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_713
timestamp 1644511149
transform 1 0 66700 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_725
timestamp 1644511149
transform 1 0 67804 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_737
timestamp 1644511149
transform 1 0 68908 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_749
timestamp 1644511149
transform 1 0 70012 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_755
timestamp 1644511149
transform 1 0 70564 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_98_757
timestamp 1644511149
transform 1 0 70748 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_769
timestamp 1644511149
transform 1 0 71852 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_781
timestamp 1644511149
transform 1 0 72956 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_793
timestamp 1644511149
transform 1 0 74060 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_805
timestamp 1644511149
transform 1 0 75164 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_811
timestamp 1644511149
transform 1 0 75716 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_98_813
timestamp 1644511149
transform 1 0 75900 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_825
timestamp 1644511149
transform 1 0 77004 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_98_837
timestamp 1644511149
transform 1 0 78108 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_98_841
timestamp 1644511149
transform 1 0 78476 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_99_3
timestamp 1644511149
transform 1 0 1380 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_15
timestamp 1644511149
transform 1 0 2484 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_27
timestamp 1644511149
transform 1 0 3588 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_39
timestamp 1644511149
transform 1 0 4692 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_99_51
timestamp 1644511149
transform 1 0 5796 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_99_55
timestamp 1644511149
transform 1 0 6164 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_99_57
timestamp 1644511149
transform 1 0 6348 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_69
timestamp 1644511149
transform 1 0 7452 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_81
timestamp 1644511149
transform 1 0 8556 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_93
timestamp 1644511149
transform 1 0 9660 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_105
timestamp 1644511149
transform 1 0 10764 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_111
timestamp 1644511149
transform 1 0 11316 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_99_113
timestamp 1644511149
transform 1 0 11500 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_125
timestamp 1644511149
transform 1 0 12604 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_137
timestamp 1644511149
transform 1 0 13708 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_149
timestamp 1644511149
transform 1 0 14812 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_161
timestamp 1644511149
transform 1 0 15916 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_167
timestamp 1644511149
transform 1 0 16468 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_99_169
timestamp 1644511149
transform 1 0 16652 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_181
timestamp 1644511149
transform 1 0 17756 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_193
timestamp 1644511149
transform 1 0 18860 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_205
timestamp 1644511149
transform 1 0 19964 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_217
timestamp 1644511149
transform 1 0 21068 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_223
timestamp 1644511149
transform 1 0 21620 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_99_225
timestamp 1644511149
transform 1 0 21804 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_237
timestamp 1644511149
transform 1 0 22908 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_249
timestamp 1644511149
transform 1 0 24012 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_261
timestamp 1644511149
transform 1 0 25116 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_273
timestamp 1644511149
transform 1 0 26220 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_279
timestamp 1644511149
transform 1 0 26772 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_99_281
timestamp 1644511149
transform 1 0 26956 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_293
timestamp 1644511149
transform 1 0 28060 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_305
timestamp 1644511149
transform 1 0 29164 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_317
timestamp 1644511149
transform 1 0 30268 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_329
timestamp 1644511149
transform 1 0 31372 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_335
timestamp 1644511149
transform 1 0 31924 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_99_337
timestamp 1644511149
transform 1 0 32108 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_349
timestamp 1644511149
transform 1 0 33212 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_361
timestamp 1644511149
transform 1 0 34316 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_373
timestamp 1644511149
transform 1 0 35420 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_385
timestamp 1644511149
transform 1 0 36524 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_391
timestamp 1644511149
transform 1 0 37076 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_99_393
timestamp 1644511149
transform 1 0 37260 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_405
timestamp 1644511149
transform 1 0 38364 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_417
timestamp 1644511149
transform 1 0 39468 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_429
timestamp 1644511149
transform 1 0 40572 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_441
timestamp 1644511149
transform 1 0 41676 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_447
timestamp 1644511149
transform 1 0 42228 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_99_449
timestamp 1644511149
transform 1 0 42412 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_461
timestamp 1644511149
transform 1 0 43516 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_473
timestamp 1644511149
transform 1 0 44620 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_485
timestamp 1644511149
transform 1 0 45724 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_497
timestamp 1644511149
transform 1 0 46828 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_503
timestamp 1644511149
transform 1 0 47380 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_99_505
timestamp 1644511149
transform 1 0 47564 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_517
timestamp 1644511149
transform 1 0 48668 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_529
timestamp 1644511149
transform 1 0 49772 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_541
timestamp 1644511149
transform 1 0 50876 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_553
timestamp 1644511149
transform 1 0 51980 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_559
timestamp 1644511149
transform 1 0 52532 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_99_561
timestamp 1644511149
transform 1 0 52716 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_573
timestamp 1644511149
transform 1 0 53820 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_585
timestamp 1644511149
transform 1 0 54924 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_597
timestamp 1644511149
transform 1 0 56028 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_609
timestamp 1644511149
transform 1 0 57132 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_615
timestamp 1644511149
transform 1 0 57684 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_99_617
timestamp 1644511149
transform 1 0 57868 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_629
timestamp 1644511149
transform 1 0 58972 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_641
timestamp 1644511149
transform 1 0 60076 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_653
timestamp 1644511149
transform 1 0 61180 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_665
timestamp 1644511149
transform 1 0 62284 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_671
timestamp 1644511149
transform 1 0 62836 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_99_673
timestamp 1644511149
transform 1 0 63020 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_685
timestamp 1644511149
transform 1 0 64124 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_697
timestamp 1644511149
transform 1 0 65228 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_709
timestamp 1644511149
transform 1 0 66332 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_721
timestamp 1644511149
transform 1 0 67436 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_727
timestamp 1644511149
transform 1 0 67988 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_99_729
timestamp 1644511149
transform 1 0 68172 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_741
timestamp 1644511149
transform 1 0 69276 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_753
timestamp 1644511149
transform 1 0 70380 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_765
timestamp 1644511149
transform 1 0 71484 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_777
timestamp 1644511149
transform 1 0 72588 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_783
timestamp 1644511149
transform 1 0 73140 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_99_785
timestamp 1644511149
transform 1 0 73324 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_797
timestamp 1644511149
transform 1 0 74428 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_809
timestamp 1644511149
transform 1 0 75532 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_99_821
timestamp 1644511149
transform 1 0 76636 0 -1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_99_829
timestamp 1644511149
transform 1 0 77372 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_99_836
timestamp 1644511149
transform 1 0 78016 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_99_841
timestamp 1644511149
transform 1 0 78476 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_100_3
timestamp 1644511149
transform 1 0 1380 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_15
timestamp 1644511149
transform 1 0 2484 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_100_27
timestamp 1644511149
transform 1 0 3588 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_100_29
timestamp 1644511149
transform 1 0 3772 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_41
timestamp 1644511149
transform 1 0 4876 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_53
timestamp 1644511149
transform 1 0 5980 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_65
timestamp 1644511149
transform 1 0 7084 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_77
timestamp 1644511149
transform 1 0 8188 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_83
timestamp 1644511149
transform 1 0 8740 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_100_85
timestamp 1644511149
transform 1 0 8924 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_97
timestamp 1644511149
transform 1 0 10028 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_109
timestamp 1644511149
transform 1 0 11132 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_121
timestamp 1644511149
transform 1 0 12236 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_133
timestamp 1644511149
transform 1 0 13340 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_139
timestamp 1644511149
transform 1 0 13892 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_100_141
timestamp 1644511149
transform 1 0 14076 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_153
timestamp 1644511149
transform 1 0 15180 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_165
timestamp 1644511149
transform 1 0 16284 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_177
timestamp 1644511149
transform 1 0 17388 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_189
timestamp 1644511149
transform 1 0 18492 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_195
timestamp 1644511149
transform 1 0 19044 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_100_197
timestamp 1644511149
transform 1 0 19228 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_209
timestamp 1644511149
transform 1 0 20332 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_221
timestamp 1644511149
transform 1 0 21436 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_233
timestamp 1644511149
transform 1 0 22540 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_245
timestamp 1644511149
transform 1 0 23644 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_251
timestamp 1644511149
transform 1 0 24196 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_100_253
timestamp 1644511149
transform 1 0 24380 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_265
timestamp 1644511149
transform 1 0 25484 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_277
timestamp 1644511149
transform 1 0 26588 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_289
timestamp 1644511149
transform 1 0 27692 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_301
timestamp 1644511149
transform 1 0 28796 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_307
timestamp 1644511149
transform 1 0 29348 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_100_309
timestamp 1644511149
transform 1 0 29532 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_321
timestamp 1644511149
transform 1 0 30636 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_333
timestamp 1644511149
transform 1 0 31740 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_345
timestamp 1644511149
transform 1 0 32844 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_357
timestamp 1644511149
transform 1 0 33948 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_363
timestamp 1644511149
transform 1 0 34500 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_100_365
timestamp 1644511149
transform 1 0 34684 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_377
timestamp 1644511149
transform 1 0 35788 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_389
timestamp 1644511149
transform 1 0 36892 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_401
timestamp 1644511149
transform 1 0 37996 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_413
timestamp 1644511149
transform 1 0 39100 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_419
timestamp 1644511149
transform 1 0 39652 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_100_421
timestamp 1644511149
transform 1 0 39836 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_433
timestamp 1644511149
transform 1 0 40940 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_445
timestamp 1644511149
transform 1 0 42044 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_457
timestamp 1644511149
transform 1 0 43148 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_469
timestamp 1644511149
transform 1 0 44252 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_475
timestamp 1644511149
transform 1 0 44804 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_100_477
timestamp 1644511149
transform 1 0 44988 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_489
timestamp 1644511149
transform 1 0 46092 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_501
timestamp 1644511149
transform 1 0 47196 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_513
timestamp 1644511149
transform 1 0 48300 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_525
timestamp 1644511149
transform 1 0 49404 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_531
timestamp 1644511149
transform 1 0 49956 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_100_533
timestamp 1644511149
transform 1 0 50140 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_545
timestamp 1644511149
transform 1 0 51244 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_557
timestamp 1644511149
transform 1 0 52348 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_569
timestamp 1644511149
transform 1 0 53452 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_581
timestamp 1644511149
transform 1 0 54556 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_587
timestamp 1644511149
transform 1 0 55108 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_100_589
timestamp 1644511149
transform 1 0 55292 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_601
timestamp 1644511149
transform 1 0 56396 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_613
timestamp 1644511149
transform 1 0 57500 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_625
timestamp 1644511149
transform 1 0 58604 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_637
timestamp 1644511149
transform 1 0 59708 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_643
timestamp 1644511149
transform 1 0 60260 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_100_645
timestamp 1644511149
transform 1 0 60444 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_657
timestamp 1644511149
transform 1 0 61548 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_669
timestamp 1644511149
transform 1 0 62652 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_681
timestamp 1644511149
transform 1 0 63756 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_693
timestamp 1644511149
transform 1 0 64860 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_699
timestamp 1644511149
transform 1 0 65412 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_100_701
timestamp 1644511149
transform 1 0 65596 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_713
timestamp 1644511149
transform 1 0 66700 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_725
timestamp 1644511149
transform 1 0 67804 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_737
timestamp 1644511149
transform 1 0 68908 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_749
timestamp 1644511149
transform 1 0 70012 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_755
timestamp 1644511149
transform 1 0 70564 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_100_757
timestamp 1644511149
transform 1 0 70748 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_769
timestamp 1644511149
transform 1 0 71852 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_781
timestamp 1644511149
transform 1 0 72956 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_793
timestamp 1644511149
transform 1 0 74060 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_805
timestamp 1644511149
transform 1 0 75164 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_811
timestamp 1644511149
transform 1 0 75716 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_100_813
timestamp 1644511149
transform 1 0 75900 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_825
timestamp 1644511149
transform 1 0 77004 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_100_837
timestamp 1644511149
transform 1 0 78108 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_100_841
timestamp 1644511149
transform 1 0 78476 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_101_3
timestamp 1644511149
transform 1 0 1380 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_15
timestamp 1644511149
transform 1 0 2484 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_27
timestamp 1644511149
transform 1 0 3588 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_39
timestamp 1644511149
transform 1 0 4692 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_101_51
timestamp 1644511149
transform 1 0 5796 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_101_55
timestamp 1644511149
transform 1 0 6164 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_101_57
timestamp 1644511149
transform 1 0 6348 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_69
timestamp 1644511149
transform 1 0 7452 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_81
timestamp 1644511149
transform 1 0 8556 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_93
timestamp 1644511149
transform 1 0 9660 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_101_105
timestamp 1644511149
transform 1 0 10764 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_111
timestamp 1644511149
transform 1 0 11316 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_101_113
timestamp 1644511149
transform 1 0 11500 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_125
timestamp 1644511149
transform 1 0 12604 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_137
timestamp 1644511149
transform 1 0 13708 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_149
timestamp 1644511149
transform 1 0 14812 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_101_161
timestamp 1644511149
transform 1 0 15916 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_167
timestamp 1644511149
transform 1 0 16468 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_101_169
timestamp 1644511149
transform 1 0 16652 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_181
timestamp 1644511149
transform 1 0 17756 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_193
timestamp 1644511149
transform 1 0 18860 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_205
timestamp 1644511149
transform 1 0 19964 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_101_217
timestamp 1644511149
transform 1 0 21068 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_223
timestamp 1644511149
transform 1 0 21620 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_101_225
timestamp 1644511149
transform 1 0 21804 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_237
timestamp 1644511149
transform 1 0 22908 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_249
timestamp 1644511149
transform 1 0 24012 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_261
timestamp 1644511149
transform 1 0 25116 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_101_273
timestamp 1644511149
transform 1 0 26220 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_279
timestamp 1644511149
transform 1 0 26772 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_101_281
timestamp 1644511149
transform 1 0 26956 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_293
timestamp 1644511149
transform 1 0 28060 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_305
timestamp 1644511149
transform 1 0 29164 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_317
timestamp 1644511149
transform 1 0 30268 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_101_329
timestamp 1644511149
transform 1 0 31372 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_335
timestamp 1644511149
transform 1 0 31924 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_101_337
timestamp 1644511149
transform 1 0 32108 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_349
timestamp 1644511149
transform 1 0 33212 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_361
timestamp 1644511149
transform 1 0 34316 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_373
timestamp 1644511149
transform 1 0 35420 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_101_385
timestamp 1644511149
transform 1 0 36524 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_391
timestamp 1644511149
transform 1 0 37076 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_101_393
timestamp 1644511149
transform 1 0 37260 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_405
timestamp 1644511149
transform 1 0 38364 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_417
timestamp 1644511149
transform 1 0 39468 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_429
timestamp 1644511149
transform 1 0 40572 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_101_441
timestamp 1644511149
transform 1 0 41676 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_447
timestamp 1644511149
transform 1 0 42228 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_101_449
timestamp 1644511149
transform 1 0 42412 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_461
timestamp 1644511149
transform 1 0 43516 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_473
timestamp 1644511149
transform 1 0 44620 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_485
timestamp 1644511149
transform 1 0 45724 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_101_497
timestamp 1644511149
transform 1 0 46828 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_503
timestamp 1644511149
transform 1 0 47380 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_101_505
timestamp 1644511149
transform 1 0 47564 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_517
timestamp 1644511149
transform 1 0 48668 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_529
timestamp 1644511149
transform 1 0 49772 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_541
timestamp 1644511149
transform 1 0 50876 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_101_553
timestamp 1644511149
transform 1 0 51980 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_559
timestamp 1644511149
transform 1 0 52532 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_101_561
timestamp 1644511149
transform 1 0 52716 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_573
timestamp 1644511149
transform 1 0 53820 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_585
timestamp 1644511149
transform 1 0 54924 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_597
timestamp 1644511149
transform 1 0 56028 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_101_609
timestamp 1644511149
transform 1 0 57132 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_615
timestamp 1644511149
transform 1 0 57684 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_101_617
timestamp 1644511149
transform 1 0 57868 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_629
timestamp 1644511149
transform 1 0 58972 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_641
timestamp 1644511149
transform 1 0 60076 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_653
timestamp 1644511149
transform 1 0 61180 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_101_665
timestamp 1644511149
transform 1 0 62284 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_671
timestamp 1644511149
transform 1 0 62836 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_101_673
timestamp 1644511149
transform 1 0 63020 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_685
timestamp 1644511149
transform 1 0 64124 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_697
timestamp 1644511149
transform 1 0 65228 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_709
timestamp 1644511149
transform 1 0 66332 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_101_721
timestamp 1644511149
transform 1 0 67436 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_727
timestamp 1644511149
transform 1 0 67988 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_101_729
timestamp 1644511149
transform 1 0 68172 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_741
timestamp 1644511149
transform 1 0 69276 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_753
timestamp 1644511149
transform 1 0 70380 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_765
timestamp 1644511149
transform 1 0 71484 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_101_777
timestamp 1644511149
transform 1 0 72588 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_783
timestamp 1644511149
transform 1 0 73140 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_101_785
timestamp 1644511149
transform 1 0 73324 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_797
timestamp 1644511149
transform 1 0 74428 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_809
timestamp 1644511149
transform 1 0 75532 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_821
timestamp 1644511149
transform 1 0 76636 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_101_833
timestamp 1644511149
transform 1 0 77740 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_839
timestamp 1644511149
transform 1 0 78292 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_101_841
timestamp 1644511149
transform 1 0 78476 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_102_3
timestamp 1644511149
transform 1 0 1380 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_15
timestamp 1644511149
transform 1 0 2484 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_102_27
timestamp 1644511149
transform 1 0 3588 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_102_29
timestamp 1644511149
transform 1 0 3772 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_41
timestamp 1644511149
transform 1 0 4876 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_53
timestamp 1644511149
transform 1 0 5980 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_65
timestamp 1644511149
transform 1 0 7084 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_102_77
timestamp 1644511149
transform 1 0 8188 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_102_83
timestamp 1644511149
transform 1 0 8740 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_102_85
timestamp 1644511149
transform 1 0 8924 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_97
timestamp 1644511149
transform 1 0 10028 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_109
timestamp 1644511149
transform 1 0 11132 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_121
timestamp 1644511149
transform 1 0 12236 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_102_133
timestamp 1644511149
transform 1 0 13340 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_102_139
timestamp 1644511149
transform 1 0 13892 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_102_141
timestamp 1644511149
transform 1 0 14076 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_153
timestamp 1644511149
transform 1 0 15180 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_165
timestamp 1644511149
transform 1 0 16284 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_177
timestamp 1644511149
transform 1 0 17388 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_102_189
timestamp 1644511149
transform 1 0 18492 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_102_195
timestamp 1644511149
transform 1 0 19044 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_102_197
timestamp 1644511149
transform 1 0 19228 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_209
timestamp 1644511149
transform 1 0 20332 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_221
timestamp 1644511149
transform 1 0 21436 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_233
timestamp 1644511149
transform 1 0 22540 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_102_245
timestamp 1644511149
transform 1 0 23644 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_102_251
timestamp 1644511149
transform 1 0 24196 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_102_253
timestamp 1644511149
transform 1 0 24380 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_265
timestamp 1644511149
transform 1 0 25484 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_277
timestamp 1644511149
transform 1 0 26588 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_289
timestamp 1644511149
transform 1 0 27692 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_102_301
timestamp 1644511149
transform 1 0 28796 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_102_307
timestamp 1644511149
transform 1 0 29348 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_102_309
timestamp 1644511149
transform 1 0 29532 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_321
timestamp 1644511149
transform 1 0 30636 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_333
timestamp 1644511149
transform 1 0 31740 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_345
timestamp 1644511149
transform 1 0 32844 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_102_357
timestamp 1644511149
transform 1 0 33948 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_102_363
timestamp 1644511149
transform 1 0 34500 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_102_365
timestamp 1644511149
transform 1 0 34684 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_377
timestamp 1644511149
transform 1 0 35788 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_389
timestamp 1644511149
transform 1 0 36892 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_401
timestamp 1644511149
transform 1 0 37996 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_102_413
timestamp 1644511149
transform 1 0 39100 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_102_419
timestamp 1644511149
transform 1 0 39652 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_102_421
timestamp 1644511149
transform 1 0 39836 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_433
timestamp 1644511149
transform 1 0 40940 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_445
timestamp 1644511149
transform 1 0 42044 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_457
timestamp 1644511149
transform 1 0 43148 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_102_469
timestamp 1644511149
transform 1 0 44252 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_102_475
timestamp 1644511149
transform 1 0 44804 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_102_477
timestamp 1644511149
transform 1 0 44988 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_489
timestamp 1644511149
transform 1 0 46092 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_501
timestamp 1644511149
transform 1 0 47196 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_513
timestamp 1644511149
transform 1 0 48300 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_102_525
timestamp 1644511149
transform 1 0 49404 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_102_531
timestamp 1644511149
transform 1 0 49956 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_102_533
timestamp 1644511149
transform 1 0 50140 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_545
timestamp 1644511149
transform 1 0 51244 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_557
timestamp 1644511149
transform 1 0 52348 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_569
timestamp 1644511149
transform 1 0 53452 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_102_581
timestamp 1644511149
transform 1 0 54556 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_102_587
timestamp 1644511149
transform 1 0 55108 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_102_589
timestamp 1644511149
transform 1 0 55292 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_601
timestamp 1644511149
transform 1 0 56396 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_613
timestamp 1644511149
transform 1 0 57500 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_625
timestamp 1644511149
transform 1 0 58604 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_102_637
timestamp 1644511149
transform 1 0 59708 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_102_643
timestamp 1644511149
transform 1 0 60260 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_102_645
timestamp 1644511149
transform 1 0 60444 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_657
timestamp 1644511149
transform 1 0 61548 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_669
timestamp 1644511149
transform 1 0 62652 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_681
timestamp 1644511149
transform 1 0 63756 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_102_693
timestamp 1644511149
transform 1 0 64860 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_102_699
timestamp 1644511149
transform 1 0 65412 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_102_701
timestamp 1644511149
transform 1 0 65596 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_713
timestamp 1644511149
transform 1 0 66700 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_725
timestamp 1644511149
transform 1 0 67804 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_737
timestamp 1644511149
transform 1 0 68908 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_102_749
timestamp 1644511149
transform 1 0 70012 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_102_755
timestamp 1644511149
transform 1 0 70564 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_102_757
timestamp 1644511149
transform 1 0 70748 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_769
timestamp 1644511149
transform 1 0 71852 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_781
timestamp 1644511149
transform 1 0 72956 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_793
timestamp 1644511149
transform 1 0 74060 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_102_805
timestamp 1644511149
transform 1 0 75164 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_102_811
timestamp 1644511149
transform 1 0 75716 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_102_813
timestamp 1644511149
transform 1 0 75900 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_825
timestamp 1644511149
transform 1 0 77004 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_102_837
timestamp 1644511149
transform 1 0 78108 0 1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_102_841
timestamp 1644511149
transform 1 0 78476 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_103_3
timestamp 1644511149
transform 1 0 1380 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_103_15
timestamp 1644511149
transform 1 0 2484 0 -1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_103_21
timestamp 1644511149
transform 1 0 3036 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_33
timestamp 1644511149
transform 1 0 4140 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_103_45
timestamp 1644511149
transform 1 0 5244 0 -1 58752
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_103_53
timestamp 1644511149
transform 1 0 5980 0 -1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_103_57
timestamp 1644511149
transform 1 0 6348 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_69
timestamp 1644511149
transform 1 0 7452 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_81
timestamp 1644511149
transform 1 0 8556 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_93
timestamp 1644511149
transform 1 0 9660 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_103_105
timestamp 1644511149
transform 1 0 10764 0 -1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_103_111
timestamp 1644511149
transform 1 0 11316 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_103_113
timestamp 1644511149
transform 1 0 11500 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_125
timestamp 1644511149
transform 1 0 12604 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_137
timestamp 1644511149
transform 1 0 13708 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_149
timestamp 1644511149
transform 1 0 14812 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_103_161
timestamp 1644511149
transform 1 0 15916 0 -1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_103_167
timestamp 1644511149
transform 1 0 16468 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_103_169
timestamp 1644511149
transform 1 0 16652 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_181
timestamp 1644511149
transform 1 0 17756 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_193
timestamp 1644511149
transform 1 0 18860 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_205
timestamp 1644511149
transform 1 0 19964 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_103_217
timestamp 1644511149
transform 1 0 21068 0 -1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_103_223
timestamp 1644511149
transform 1 0 21620 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_103_225
timestamp 1644511149
transform 1 0 21804 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_237
timestamp 1644511149
transform 1 0 22908 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_249
timestamp 1644511149
transform 1 0 24012 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_261
timestamp 1644511149
transform 1 0 25116 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_103_273
timestamp 1644511149
transform 1 0 26220 0 -1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_103_279
timestamp 1644511149
transform 1 0 26772 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_103_281
timestamp 1644511149
transform 1 0 26956 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_293
timestamp 1644511149
transform 1 0 28060 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_305
timestamp 1644511149
transform 1 0 29164 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_317
timestamp 1644511149
transform 1 0 30268 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_103_329
timestamp 1644511149
transform 1 0 31372 0 -1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_103_335
timestamp 1644511149
transform 1 0 31924 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_103_337
timestamp 1644511149
transform 1 0 32108 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_349
timestamp 1644511149
transform 1 0 33212 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_361
timestamp 1644511149
transform 1 0 34316 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_373
timestamp 1644511149
transform 1 0 35420 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_103_385
timestamp 1644511149
transform 1 0 36524 0 -1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_103_391
timestamp 1644511149
transform 1 0 37076 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_103_393
timestamp 1644511149
transform 1 0 37260 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_405
timestamp 1644511149
transform 1 0 38364 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_417
timestamp 1644511149
transform 1 0 39468 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_429
timestamp 1644511149
transform 1 0 40572 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_103_441
timestamp 1644511149
transform 1 0 41676 0 -1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_103_447
timestamp 1644511149
transform 1 0 42228 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_103_449
timestamp 1644511149
transform 1 0 42412 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_461
timestamp 1644511149
transform 1 0 43516 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_473
timestamp 1644511149
transform 1 0 44620 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_485
timestamp 1644511149
transform 1 0 45724 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_103_497
timestamp 1644511149
transform 1 0 46828 0 -1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_103_503
timestamp 1644511149
transform 1 0 47380 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_103_505
timestamp 1644511149
transform 1 0 47564 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_517
timestamp 1644511149
transform 1 0 48668 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_529
timestamp 1644511149
transform 1 0 49772 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_541
timestamp 1644511149
transform 1 0 50876 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_103_553
timestamp 1644511149
transform 1 0 51980 0 -1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_103_559
timestamp 1644511149
transform 1 0 52532 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_103_561
timestamp 1644511149
transform 1 0 52716 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_573
timestamp 1644511149
transform 1 0 53820 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_585
timestamp 1644511149
transform 1 0 54924 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_597
timestamp 1644511149
transform 1 0 56028 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_103_609
timestamp 1644511149
transform 1 0 57132 0 -1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_103_615
timestamp 1644511149
transform 1 0 57684 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_103_617
timestamp 1644511149
transform 1 0 57868 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_629
timestamp 1644511149
transform 1 0 58972 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_641
timestamp 1644511149
transform 1 0 60076 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_653
timestamp 1644511149
transform 1 0 61180 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_103_665
timestamp 1644511149
transform 1 0 62284 0 -1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_103_671
timestamp 1644511149
transform 1 0 62836 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_103_673
timestamp 1644511149
transform 1 0 63020 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_685
timestamp 1644511149
transform 1 0 64124 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_697
timestamp 1644511149
transform 1 0 65228 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_709
timestamp 1644511149
transform 1 0 66332 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_103_721
timestamp 1644511149
transform 1 0 67436 0 -1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_103_727
timestamp 1644511149
transform 1 0 67988 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_103_729
timestamp 1644511149
transform 1 0 68172 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_741
timestamp 1644511149
transform 1 0 69276 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_753
timestamp 1644511149
transform 1 0 70380 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_765
timestamp 1644511149
transform 1 0 71484 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_103_777
timestamp 1644511149
transform 1 0 72588 0 -1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_103_783
timestamp 1644511149
transform 1 0 73140 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_103_785
timestamp 1644511149
transform 1 0 73324 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_797
timestamp 1644511149
transform 1 0 74428 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_809
timestamp 1644511149
transform 1 0 75532 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_821
timestamp 1644511149
transform 1 0 76636 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_103_833
timestamp 1644511149
transform 1 0 77740 0 -1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_103_839
timestamp 1644511149
transform 1 0 78292 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_103_841
timestamp 1644511149
transform 1 0 78476 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_104_7
timestamp 1644511149
transform 1 0 1748 0 1 58752
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_104_15
timestamp 1644511149
transform 1 0 2484 0 1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_104_22
timestamp 1644511149
transform 1 0 3128 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_104_29
timestamp 1644511149
transform 1 0 3772 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_41
timestamp 1644511149
transform 1 0 4876 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_53
timestamp 1644511149
transform 1 0 5980 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_65
timestamp 1644511149
transform 1 0 7084 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_104_77
timestamp 1644511149
transform 1 0 8188 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_104_83
timestamp 1644511149
transform 1 0 8740 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_104_85
timestamp 1644511149
transform 1 0 8924 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_97
timestamp 1644511149
transform 1 0 10028 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_109
timestamp 1644511149
transform 1 0 11132 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_121
timestamp 1644511149
transform 1 0 12236 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_104_133
timestamp 1644511149
transform 1 0 13340 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_104_139
timestamp 1644511149
transform 1 0 13892 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_104_141
timestamp 1644511149
transform 1 0 14076 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_153
timestamp 1644511149
transform 1 0 15180 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_165
timestamp 1644511149
transform 1 0 16284 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_177
timestamp 1644511149
transform 1 0 17388 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_104_189
timestamp 1644511149
transform 1 0 18492 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_104_195
timestamp 1644511149
transform 1 0 19044 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_104_197
timestamp 1644511149
transform 1 0 19228 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_209
timestamp 1644511149
transform 1 0 20332 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_221
timestamp 1644511149
transform 1 0 21436 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_233
timestamp 1644511149
transform 1 0 22540 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_104_245
timestamp 1644511149
transform 1 0 23644 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_104_251
timestamp 1644511149
transform 1 0 24196 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_104_253
timestamp 1644511149
transform 1 0 24380 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_265
timestamp 1644511149
transform 1 0 25484 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_277
timestamp 1644511149
transform 1 0 26588 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_289
timestamp 1644511149
transform 1 0 27692 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_104_301
timestamp 1644511149
transform 1 0 28796 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_104_307
timestamp 1644511149
transform 1 0 29348 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_104_309
timestamp 1644511149
transform 1 0 29532 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_321
timestamp 1644511149
transform 1 0 30636 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_333
timestamp 1644511149
transform 1 0 31740 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_345
timestamp 1644511149
transform 1 0 32844 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_104_357
timestamp 1644511149
transform 1 0 33948 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_104_363
timestamp 1644511149
transform 1 0 34500 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_104_365
timestamp 1644511149
transform 1 0 34684 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_377
timestamp 1644511149
transform 1 0 35788 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_389
timestamp 1644511149
transform 1 0 36892 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_401
timestamp 1644511149
transform 1 0 37996 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_104_413
timestamp 1644511149
transform 1 0 39100 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_104_419
timestamp 1644511149
transform 1 0 39652 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_104_427
timestamp 1644511149
transform 1 0 40388 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_439
timestamp 1644511149
transform 1 0 41492 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_451
timestamp 1644511149
transform 1 0 42596 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_463
timestamp 1644511149
transform 1 0 43700 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_104_475
timestamp 1644511149
transform 1 0 44804 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_104_477
timestamp 1644511149
transform 1 0 44988 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_489
timestamp 1644511149
transform 1 0 46092 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_501
timestamp 1644511149
transform 1 0 47196 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_513
timestamp 1644511149
transform 1 0 48300 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_104_525
timestamp 1644511149
transform 1 0 49404 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_104_531
timestamp 1644511149
transform 1 0 49956 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_104_533
timestamp 1644511149
transform 1 0 50140 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_545
timestamp 1644511149
transform 1 0 51244 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_557
timestamp 1644511149
transform 1 0 52348 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_569
timestamp 1644511149
transform 1 0 53452 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_104_581
timestamp 1644511149
transform 1 0 54556 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_104_587
timestamp 1644511149
transform 1 0 55108 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_104_589
timestamp 1644511149
transform 1 0 55292 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_601
timestamp 1644511149
transform 1 0 56396 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_613
timestamp 1644511149
transform 1 0 57500 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_625
timestamp 1644511149
transform 1 0 58604 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_104_637
timestamp 1644511149
transform 1 0 59708 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_104_643
timestamp 1644511149
transform 1 0 60260 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_104_645
timestamp 1644511149
transform 1 0 60444 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_657
timestamp 1644511149
transform 1 0 61548 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_669
timestamp 1644511149
transform 1 0 62652 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_681
timestamp 1644511149
transform 1 0 63756 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_104_693
timestamp 1644511149
transform 1 0 64860 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_104_699
timestamp 1644511149
transform 1 0 65412 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_104_701
timestamp 1644511149
transform 1 0 65596 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_713
timestamp 1644511149
transform 1 0 66700 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_725
timestamp 1644511149
transform 1 0 67804 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_737
timestamp 1644511149
transform 1 0 68908 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_104_749
timestamp 1644511149
transform 1 0 70012 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_104_755
timestamp 1644511149
transform 1 0 70564 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_104_757
timestamp 1644511149
transform 1 0 70748 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_769
timestamp 1644511149
transform 1 0 71852 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_781
timestamp 1644511149
transform 1 0 72956 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_793
timestamp 1644511149
transform 1 0 74060 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_104_805
timestamp 1644511149
transform 1 0 75164 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_104_811
timestamp 1644511149
transform 1 0 75716 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_104_813
timestamp 1644511149
transform 1 0 75900 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_825
timestamp 1644511149
transform 1 0 77004 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_104_837
timestamp 1644511149
transform 1 0 78108 0 1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_104_841
timestamp 1644511149
transform 1 0 78476 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_105_3
timestamp 1644511149
transform 1 0 1380 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_15
timestamp 1644511149
transform 1 0 2484 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_27
timestamp 1644511149
transform 1 0 3588 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_39
timestamp 1644511149
transform 1 0 4692 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_105_51
timestamp 1644511149
transform 1 0 5796 0 -1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_105_55
timestamp 1644511149
transform 1 0 6164 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_105_57
timestamp 1644511149
transform 1 0 6348 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_69
timestamp 1644511149
transform 1 0 7452 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_81
timestamp 1644511149
transform 1 0 8556 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_93
timestamp 1644511149
transform 1 0 9660 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_105_105
timestamp 1644511149
transform 1 0 10764 0 -1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_105_111
timestamp 1644511149
transform 1 0 11316 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_105_113
timestamp 1644511149
transform 1 0 11500 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_125
timestamp 1644511149
transform 1 0 12604 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_137
timestamp 1644511149
transform 1 0 13708 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_149
timestamp 1644511149
transform 1 0 14812 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_105_161
timestamp 1644511149
transform 1 0 15916 0 -1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_105_167
timestamp 1644511149
transform 1 0 16468 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_105_169
timestamp 1644511149
transform 1 0 16652 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_181
timestamp 1644511149
transform 1 0 17756 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_193
timestamp 1644511149
transform 1 0 18860 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_205
timestamp 1644511149
transform 1 0 19964 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_105_217
timestamp 1644511149
transform 1 0 21068 0 -1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_105_223
timestamp 1644511149
transform 1 0 21620 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_105_225
timestamp 1644511149
transform 1 0 21804 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_237
timestamp 1644511149
transform 1 0 22908 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_249
timestamp 1644511149
transform 1 0 24012 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_261
timestamp 1644511149
transform 1 0 25116 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_105_273
timestamp 1644511149
transform 1 0 26220 0 -1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_105_279
timestamp 1644511149
transform 1 0 26772 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_105_281
timestamp 1644511149
transform 1 0 26956 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_293
timestamp 1644511149
transform 1 0 28060 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_305
timestamp 1644511149
transform 1 0 29164 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_317
timestamp 1644511149
transform 1 0 30268 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_105_329
timestamp 1644511149
transform 1 0 31372 0 -1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_105_335
timestamp 1644511149
transform 1 0 31924 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_105_337
timestamp 1644511149
transform 1 0 32108 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_349
timestamp 1644511149
transform 1 0 33212 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_361
timestamp 1644511149
transform 1 0 34316 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_373
timestamp 1644511149
transform 1 0 35420 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_105_385
timestamp 1644511149
transform 1 0 36524 0 -1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_105_391
timestamp 1644511149
transform 1 0 37076 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_105_393
timestamp 1644511149
transform 1 0 37260 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_105_405
timestamp 1644511149
transform 1 0 38364 0 -1 59840
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_105_409
timestamp 1644511149
transform 1 0 38732 0 -1 59840
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_105_417
timestamp 1644511149
transform 1 0 39468 0 -1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_105_430
timestamp 1644511149
transform 1 0 40664 0 -1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_105_438
timestamp 1644511149
transform 1 0 41400 0 -1 59840
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_105_446
timestamp 1644511149
transform 1 0 42136 0 -1 59840
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_105_449
timestamp 1644511149
transform 1 0 42412 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_461
timestamp 1644511149
transform 1 0 43516 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_473
timestamp 1644511149
transform 1 0 44620 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_485
timestamp 1644511149
transform 1 0 45724 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_105_497
timestamp 1644511149
transform 1 0 46828 0 -1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_105_503
timestamp 1644511149
transform 1 0 47380 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_105_505
timestamp 1644511149
transform 1 0 47564 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_517
timestamp 1644511149
transform 1 0 48668 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_529
timestamp 1644511149
transform 1 0 49772 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_541
timestamp 1644511149
transform 1 0 50876 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_105_553
timestamp 1644511149
transform 1 0 51980 0 -1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_105_559
timestamp 1644511149
transform 1 0 52532 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_105_561
timestamp 1644511149
transform 1 0 52716 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_573
timestamp 1644511149
transform 1 0 53820 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_585
timestamp 1644511149
transform 1 0 54924 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_597
timestamp 1644511149
transform 1 0 56028 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_105_609
timestamp 1644511149
transform 1 0 57132 0 -1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_105_615
timestamp 1644511149
transform 1 0 57684 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_105_617
timestamp 1644511149
transform 1 0 57868 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_629
timestamp 1644511149
transform 1 0 58972 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_641
timestamp 1644511149
transform 1 0 60076 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_653
timestamp 1644511149
transform 1 0 61180 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_105_665
timestamp 1644511149
transform 1 0 62284 0 -1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_105_671
timestamp 1644511149
transform 1 0 62836 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_105_673
timestamp 1644511149
transform 1 0 63020 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_685
timestamp 1644511149
transform 1 0 64124 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_697
timestamp 1644511149
transform 1 0 65228 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_709
timestamp 1644511149
transform 1 0 66332 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_105_721
timestamp 1644511149
transform 1 0 67436 0 -1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_105_727
timestamp 1644511149
transform 1 0 67988 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_105_729
timestamp 1644511149
transform 1 0 68172 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_741
timestamp 1644511149
transform 1 0 69276 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_753
timestamp 1644511149
transform 1 0 70380 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_765
timestamp 1644511149
transform 1 0 71484 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_105_777
timestamp 1644511149
transform 1 0 72588 0 -1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_105_783
timestamp 1644511149
transform 1 0 73140 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_105_785
timestamp 1644511149
transform 1 0 73324 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_105_797
timestamp 1644511149
transform 1 0 74428 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_105_801
timestamp 1644511149
transform 1 0 74796 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_813
timestamp 1644511149
transform 1 0 75900 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_105_825
timestamp 1644511149
transform 1 0 77004 0 -1 59840
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_105_836
timestamp 1644511149
transform 1 0 78016 0 -1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_105_841
timestamp 1644511149
transform 1 0 78476 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_106_3
timestamp 1644511149
transform 1 0 1380 0 1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_106_11
timestamp 1644511149
transform 1 0 2116 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_106_23
timestamp 1644511149
transform 1 0 3220 0 1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_106_27
timestamp 1644511149
transform 1 0 3588 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_106_29
timestamp 1644511149
transform 1 0 3772 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_41
timestamp 1644511149
transform 1 0 4876 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_53
timestamp 1644511149
transform 1 0 5980 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_65
timestamp 1644511149
transform 1 0 7084 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_106_77
timestamp 1644511149
transform 1 0 8188 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_106_83
timestamp 1644511149
transform 1 0 8740 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_106_85
timestamp 1644511149
transform 1 0 8924 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_97
timestamp 1644511149
transform 1 0 10028 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_109
timestamp 1644511149
transform 1 0 11132 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_121
timestamp 1644511149
transform 1 0 12236 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_106_133
timestamp 1644511149
transform 1 0 13340 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_106_139
timestamp 1644511149
transform 1 0 13892 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_106_141
timestamp 1644511149
transform 1 0 14076 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_153
timestamp 1644511149
transform 1 0 15180 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_165
timestamp 1644511149
transform 1 0 16284 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_177
timestamp 1644511149
transform 1 0 17388 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_106_189
timestamp 1644511149
transform 1 0 18492 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_106_195
timestamp 1644511149
transform 1 0 19044 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_106_203
timestamp 1644511149
transform 1 0 19780 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_215
timestamp 1644511149
transform 1 0 20884 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_227
timestamp 1644511149
transform 1 0 21988 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_239
timestamp 1644511149
transform 1 0 23092 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_106_251
timestamp 1644511149
transform 1 0 24196 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_106_253
timestamp 1644511149
transform 1 0 24380 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_265
timestamp 1644511149
transform 1 0 25484 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_277
timestamp 1644511149
transform 1 0 26588 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_289
timestamp 1644511149
transform 1 0 27692 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_106_301
timestamp 1644511149
transform 1 0 28796 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_106_307
timestamp 1644511149
transform 1 0 29348 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_106_309
timestamp 1644511149
transform 1 0 29532 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_321
timestamp 1644511149
transform 1 0 30636 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_333
timestamp 1644511149
transform 1 0 31740 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_345
timestamp 1644511149
transform 1 0 32844 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_106_357
timestamp 1644511149
transform 1 0 33948 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_106_363
timestamp 1644511149
transform 1 0 34500 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_106_365
timestamp 1644511149
transform 1 0 34684 0 1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_106_375
timestamp 1644511149
transform 1 0 35604 0 1 59840
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_106_379
timestamp 1644511149
transform 1 0 35972 0 1 59840
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_106_387
timestamp 1644511149
transform 1 0 36708 0 1 59840
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_106_395
timestamp 1644511149
transform 1 0 37444 0 1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_106_400
timestamp 1644511149
transform 1 0 37904 0 1 59840
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_106_406
timestamp 1644511149
transform 1 0 38456 0 1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_106_416
timestamp 1644511149
transform 1 0 39376 0 1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_106_430
timestamp 1644511149
transform 1 0 40664 0 1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_106_440
timestamp 1644511149
transform 1 0 41584 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_452
timestamp 1644511149
transform 1 0 42688 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_464
timestamp 1644511149
transform 1 0 43792 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_477
timestamp 1644511149
transform 1 0 44988 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_489
timestamp 1644511149
transform 1 0 46092 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_501
timestamp 1644511149
transform 1 0 47196 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_513
timestamp 1644511149
transform 1 0 48300 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_106_525
timestamp 1644511149
transform 1 0 49404 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_106_531
timestamp 1644511149
transform 1 0 49956 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_106_533
timestamp 1644511149
transform 1 0 50140 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_545
timestamp 1644511149
transform 1 0 51244 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_557
timestamp 1644511149
transform 1 0 52348 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_569
timestamp 1644511149
transform 1 0 53452 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_106_581
timestamp 1644511149
transform 1 0 54556 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_106_587
timestamp 1644511149
transform 1 0 55108 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_106_589
timestamp 1644511149
transform 1 0 55292 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_601
timestamp 1644511149
transform 1 0 56396 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_613
timestamp 1644511149
transform 1 0 57500 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_625
timestamp 1644511149
transform 1 0 58604 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_106_637
timestamp 1644511149
transform 1 0 59708 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_106_643
timestamp 1644511149
transform 1 0 60260 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_106_645
timestamp 1644511149
transform 1 0 60444 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_657
timestamp 1644511149
transform 1 0 61548 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_106_669
timestamp 1644511149
transform 1 0 62652 0 1 59840
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_106_677
timestamp 1644511149
transform 1 0 63388 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_106_689
timestamp 1644511149
transform 1 0 64492 0 1 59840
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_106_697
timestamp 1644511149
transform 1 0 65228 0 1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_106_701
timestamp 1644511149
transform 1 0 65596 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_713
timestamp 1644511149
transform 1 0 66700 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_725
timestamp 1644511149
transform 1 0 67804 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_737
timestamp 1644511149
transform 1 0 68908 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_106_749
timestamp 1644511149
transform 1 0 70012 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_106_755
timestamp 1644511149
transform 1 0 70564 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_106_757
timestamp 1644511149
transform 1 0 70748 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_769
timestamp 1644511149
transform 1 0 71852 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_781
timestamp 1644511149
transform 1 0 72956 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_793
timestamp 1644511149
transform 1 0 74060 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_106_805
timestamp 1644511149
transform 1 0 75164 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_106_811
timestamp 1644511149
transform 1 0 75716 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_106_813
timestamp 1644511149
transform 1 0 75900 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_106_825
timestamp 1644511149
transform 1 0 77004 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_106_831
timestamp 1644511149
transform 1 0 77556 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_106_838
timestamp 1644511149
transform 1 0 78200 0 1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_107_3
timestamp 1644511149
transform 1 0 1380 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_15
timestamp 1644511149
transform 1 0 2484 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_27
timestamp 1644511149
transform 1 0 3588 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_39
timestamp 1644511149
transform 1 0 4692 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_107_51
timestamp 1644511149
transform 1 0 5796 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_107_55
timestamp 1644511149
transform 1 0 6164 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_107_57
timestamp 1644511149
transform 1 0 6348 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_69
timestamp 1644511149
transform 1 0 7452 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_81
timestamp 1644511149
transform 1 0 8556 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_93
timestamp 1644511149
transform 1 0 9660 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_107_105
timestamp 1644511149
transform 1 0 10764 0 -1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_107_111
timestamp 1644511149
transform 1 0 11316 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_107_113
timestamp 1644511149
transform 1 0 11500 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_125
timestamp 1644511149
transform 1 0 12604 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_137
timestamp 1644511149
transform 1 0 13708 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_149
timestamp 1644511149
transform 1 0 14812 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_107_161
timestamp 1644511149
transform 1 0 15916 0 -1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_107_167
timestamp 1644511149
transform 1 0 16468 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_107_169
timestamp 1644511149
transform 1 0 16652 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_181
timestamp 1644511149
transform 1 0 17756 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_193
timestamp 1644511149
transform 1 0 18860 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_205
timestamp 1644511149
transform 1 0 19964 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_107_217
timestamp 1644511149
transform 1 0 21068 0 -1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_107_223
timestamp 1644511149
transform 1 0 21620 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_107_225
timestamp 1644511149
transform 1 0 21804 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_237
timestamp 1644511149
transform 1 0 22908 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_249
timestamp 1644511149
transform 1 0 24012 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_261
timestamp 1644511149
transform 1 0 25116 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_107_273
timestamp 1644511149
transform 1 0 26220 0 -1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_107_279
timestamp 1644511149
transform 1 0 26772 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_107_281
timestamp 1644511149
transform 1 0 26956 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_293
timestamp 1644511149
transform 1 0 28060 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_305
timestamp 1644511149
transform 1 0 29164 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_317
timestamp 1644511149
transform 1 0 30268 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_107_329
timestamp 1644511149
transform 1 0 31372 0 -1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_107_335
timestamp 1644511149
transform 1 0 31924 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_107_337
timestamp 1644511149
transform 1 0 32108 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_349
timestamp 1644511149
transform 1 0 33212 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_361
timestamp 1644511149
transform 1 0 34316 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_373
timestamp 1644511149
transform 1 0 35420 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_107_385
timestamp 1644511149
transform 1 0 36524 0 -1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_107_391
timestamp 1644511149
transform 1 0 37076 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_107_393
timestamp 1644511149
transform 1 0 37260 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_107_405
timestamp 1644511149
transform 1 0 38364 0 -1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_107_417
timestamp 1644511149
transform 1 0 39468 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_107_427
timestamp 1644511149
transform 1 0 40388 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_107_437
timestamp 1644511149
transform 1 0 41308 0 -1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_107_445
timestamp 1644511149
transform 1 0 42044 0 -1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_107_449
timestamp 1644511149
transform 1 0 42412 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_461
timestamp 1644511149
transform 1 0 43516 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_473
timestamp 1644511149
transform 1 0 44620 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_485
timestamp 1644511149
transform 1 0 45724 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_107_497
timestamp 1644511149
transform 1 0 46828 0 -1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_107_503
timestamp 1644511149
transform 1 0 47380 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_107_505
timestamp 1644511149
transform 1 0 47564 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_517
timestamp 1644511149
transform 1 0 48668 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_529
timestamp 1644511149
transform 1 0 49772 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_541
timestamp 1644511149
transform 1 0 50876 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_107_553
timestamp 1644511149
transform 1 0 51980 0 -1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_107_559
timestamp 1644511149
transform 1 0 52532 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_107_561
timestamp 1644511149
transform 1 0 52716 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_573
timestamp 1644511149
transform 1 0 53820 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_585
timestamp 1644511149
transform 1 0 54924 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_597
timestamp 1644511149
transform 1 0 56028 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_107_609
timestamp 1644511149
transform 1 0 57132 0 -1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_107_615
timestamp 1644511149
transform 1 0 57684 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_107_617
timestamp 1644511149
transform 1 0 57868 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_629
timestamp 1644511149
transform 1 0 58972 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_641
timestamp 1644511149
transform 1 0 60076 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_653
timestamp 1644511149
transform 1 0 61180 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_107_665
timestamp 1644511149
transform 1 0 62284 0 -1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_107_671
timestamp 1644511149
transform 1 0 62836 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_107_673
timestamp 1644511149
transform 1 0 63020 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_685
timestamp 1644511149
transform 1 0 64124 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_697
timestamp 1644511149
transform 1 0 65228 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_709
timestamp 1644511149
transform 1 0 66332 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_107_721
timestamp 1644511149
transform 1 0 67436 0 -1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_107_727
timestamp 1644511149
transform 1 0 67988 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_107_729
timestamp 1644511149
transform 1 0 68172 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_741
timestamp 1644511149
transform 1 0 69276 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_753
timestamp 1644511149
transform 1 0 70380 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_765
timestamp 1644511149
transform 1 0 71484 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_107_777
timestamp 1644511149
transform 1 0 72588 0 -1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_107_783
timestamp 1644511149
transform 1 0 73140 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_107_785
timestamp 1644511149
transform 1 0 73324 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_797
timestamp 1644511149
transform 1 0 74428 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_809
timestamp 1644511149
transform 1 0 75532 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_821
timestamp 1644511149
transform 1 0 76636 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_107_833
timestamp 1644511149
transform 1 0 77740 0 -1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_107_839
timestamp 1644511149
transform 1 0 78292 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_107_841
timestamp 1644511149
transform 1 0 78476 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_108_3
timestamp 1644511149
transform 1 0 1380 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_15
timestamp 1644511149
transform 1 0 2484 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_108_27
timestamp 1644511149
transform 1 0 3588 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_108_29
timestamp 1644511149
transform 1 0 3772 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_41
timestamp 1644511149
transform 1 0 4876 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_53
timestamp 1644511149
transform 1 0 5980 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_65
timestamp 1644511149
transform 1 0 7084 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_108_77
timestamp 1644511149
transform 1 0 8188 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_108_83
timestamp 1644511149
transform 1 0 8740 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_108_85
timestamp 1644511149
transform 1 0 8924 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_97
timestamp 1644511149
transform 1 0 10028 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_109
timestamp 1644511149
transform 1 0 11132 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_121
timestamp 1644511149
transform 1 0 12236 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_108_133
timestamp 1644511149
transform 1 0 13340 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_108_139
timestamp 1644511149
transform 1 0 13892 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_108_141
timestamp 1644511149
transform 1 0 14076 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_153
timestamp 1644511149
transform 1 0 15180 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_165
timestamp 1644511149
transform 1 0 16284 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_177
timestamp 1644511149
transform 1 0 17388 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_108_189
timestamp 1644511149
transform 1 0 18492 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_108_195
timestamp 1644511149
transform 1 0 19044 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_108_197
timestamp 1644511149
transform 1 0 19228 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_209
timestamp 1644511149
transform 1 0 20332 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_221
timestamp 1644511149
transform 1 0 21436 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_233
timestamp 1644511149
transform 1 0 22540 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_108_245
timestamp 1644511149
transform 1 0 23644 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_108_251
timestamp 1644511149
transform 1 0 24196 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_108_253
timestamp 1644511149
transform 1 0 24380 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_265
timestamp 1644511149
transform 1 0 25484 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_277
timestamp 1644511149
transform 1 0 26588 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_289
timestamp 1644511149
transform 1 0 27692 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_108_301
timestamp 1644511149
transform 1 0 28796 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_108_307
timestamp 1644511149
transform 1 0 29348 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_108_309
timestamp 1644511149
transform 1 0 29532 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_321
timestamp 1644511149
transform 1 0 30636 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_333
timestamp 1644511149
transform 1 0 31740 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_345
timestamp 1644511149
transform 1 0 32844 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_108_357
timestamp 1644511149
transform 1 0 33948 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_108_363
timestamp 1644511149
transform 1 0 34500 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_108_365
timestamp 1644511149
transform 1 0 34684 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_377
timestamp 1644511149
transform 1 0 35788 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_389
timestamp 1644511149
transform 1 0 36892 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_401
timestamp 1644511149
transform 1 0 37996 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_108_413
timestamp 1644511149
transform 1 0 39100 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_108_419
timestamp 1644511149
transform 1 0 39652 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_108_427
timestamp 1644511149
transform 1 0 40388 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_439
timestamp 1644511149
transform 1 0 41492 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_451
timestamp 1644511149
transform 1 0 42596 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_463
timestamp 1644511149
transform 1 0 43700 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_108_475
timestamp 1644511149
transform 1 0 44804 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_108_477
timestamp 1644511149
transform 1 0 44988 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_489
timestamp 1644511149
transform 1 0 46092 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_501
timestamp 1644511149
transform 1 0 47196 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_513
timestamp 1644511149
transform 1 0 48300 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_108_525
timestamp 1644511149
transform 1 0 49404 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_108_531
timestamp 1644511149
transform 1 0 49956 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_108_533
timestamp 1644511149
transform 1 0 50140 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_545
timestamp 1644511149
transform 1 0 51244 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_557
timestamp 1644511149
transform 1 0 52348 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_569
timestamp 1644511149
transform 1 0 53452 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_108_581
timestamp 1644511149
transform 1 0 54556 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_108_587
timestamp 1644511149
transform 1 0 55108 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_108_589
timestamp 1644511149
transform 1 0 55292 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_601
timestamp 1644511149
transform 1 0 56396 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_613
timestamp 1644511149
transform 1 0 57500 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_625
timestamp 1644511149
transform 1 0 58604 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_108_637
timestamp 1644511149
transform 1 0 59708 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_108_643
timestamp 1644511149
transform 1 0 60260 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_108_645
timestamp 1644511149
transform 1 0 60444 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_657
timestamp 1644511149
transform 1 0 61548 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_669
timestamp 1644511149
transform 1 0 62652 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_681
timestamp 1644511149
transform 1 0 63756 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_108_693
timestamp 1644511149
transform 1 0 64860 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_108_699
timestamp 1644511149
transform 1 0 65412 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_108_701
timestamp 1644511149
transform 1 0 65596 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_713
timestamp 1644511149
transform 1 0 66700 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_725
timestamp 1644511149
transform 1 0 67804 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_737
timestamp 1644511149
transform 1 0 68908 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_108_749
timestamp 1644511149
transform 1 0 70012 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_108_755
timestamp 1644511149
transform 1 0 70564 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_108_757
timestamp 1644511149
transform 1 0 70748 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_769
timestamp 1644511149
transform 1 0 71852 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_781
timestamp 1644511149
transform 1 0 72956 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_793
timestamp 1644511149
transform 1 0 74060 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_108_805
timestamp 1644511149
transform 1 0 75164 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_108_811
timestamp 1644511149
transform 1 0 75716 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_108_813
timestamp 1644511149
transform 1 0 75900 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_825
timestamp 1644511149
transform 1 0 77004 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_108_837
timestamp 1644511149
transform 1 0 78108 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_108_841
timestamp 1644511149
transform 1 0 78476 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_109_3
timestamp 1644511149
transform 1 0 1380 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_15
timestamp 1644511149
transform 1 0 2484 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_27
timestamp 1644511149
transform 1 0 3588 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_39
timestamp 1644511149
transform 1 0 4692 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_109_51
timestamp 1644511149
transform 1 0 5796 0 -1 62016
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_109_55
timestamp 1644511149
transform 1 0 6164 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_109_57
timestamp 1644511149
transform 1 0 6348 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_69
timestamp 1644511149
transform 1 0 7452 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_81
timestamp 1644511149
transform 1 0 8556 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_93
timestamp 1644511149
transform 1 0 9660 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_109_105
timestamp 1644511149
transform 1 0 10764 0 -1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_109_111
timestamp 1644511149
transform 1 0 11316 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_109_113
timestamp 1644511149
transform 1 0 11500 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_125
timestamp 1644511149
transform 1 0 12604 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_137
timestamp 1644511149
transform 1 0 13708 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_149
timestamp 1644511149
transform 1 0 14812 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_109_161
timestamp 1644511149
transform 1 0 15916 0 -1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_109_167
timestamp 1644511149
transform 1 0 16468 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_109_169
timestamp 1644511149
transform 1 0 16652 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_181
timestamp 1644511149
transform 1 0 17756 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_193
timestamp 1644511149
transform 1 0 18860 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_205
timestamp 1644511149
transform 1 0 19964 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_109_217
timestamp 1644511149
transform 1 0 21068 0 -1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_109_223
timestamp 1644511149
transform 1 0 21620 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_109_225
timestamp 1644511149
transform 1 0 21804 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_237
timestamp 1644511149
transform 1 0 22908 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_249
timestamp 1644511149
transform 1 0 24012 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_261
timestamp 1644511149
transform 1 0 25116 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_109_273
timestamp 1644511149
transform 1 0 26220 0 -1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_109_279
timestamp 1644511149
transform 1 0 26772 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_109_281
timestamp 1644511149
transform 1 0 26956 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_293
timestamp 1644511149
transform 1 0 28060 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_305
timestamp 1644511149
transform 1 0 29164 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_317
timestamp 1644511149
transform 1 0 30268 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_109_329
timestamp 1644511149
transform 1 0 31372 0 -1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_109_335
timestamp 1644511149
transform 1 0 31924 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_109_337
timestamp 1644511149
transform 1 0 32108 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_349
timestamp 1644511149
transform 1 0 33212 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_361
timestamp 1644511149
transform 1 0 34316 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_373
timestamp 1644511149
transform 1 0 35420 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_109_385
timestamp 1644511149
transform 1 0 36524 0 -1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_109_391
timestamp 1644511149
transform 1 0 37076 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_109_393
timestamp 1644511149
transform 1 0 37260 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_405
timestamp 1644511149
transform 1 0 38364 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_417
timestamp 1644511149
transform 1 0 39468 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_429
timestamp 1644511149
transform 1 0 40572 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_109_441
timestamp 1644511149
transform 1 0 41676 0 -1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_109_447
timestamp 1644511149
transform 1 0 42228 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_109_449
timestamp 1644511149
transform 1 0 42412 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_461
timestamp 1644511149
transform 1 0 43516 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_473
timestamp 1644511149
transform 1 0 44620 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_485
timestamp 1644511149
transform 1 0 45724 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_109_497
timestamp 1644511149
transform 1 0 46828 0 -1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_109_503
timestamp 1644511149
transform 1 0 47380 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_109_505
timestamp 1644511149
transform 1 0 47564 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_517
timestamp 1644511149
transform 1 0 48668 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_529
timestamp 1644511149
transform 1 0 49772 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_541
timestamp 1644511149
transform 1 0 50876 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_109_553
timestamp 1644511149
transform 1 0 51980 0 -1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_109_559
timestamp 1644511149
transform 1 0 52532 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_109_561
timestamp 1644511149
transform 1 0 52716 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_573
timestamp 1644511149
transform 1 0 53820 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_585
timestamp 1644511149
transform 1 0 54924 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_597
timestamp 1644511149
transform 1 0 56028 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_109_609
timestamp 1644511149
transform 1 0 57132 0 -1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_109_615
timestamp 1644511149
transform 1 0 57684 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_109_617
timestamp 1644511149
transform 1 0 57868 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_629
timestamp 1644511149
transform 1 0 58972 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_641
timestamp 1644511149
transform 1 0 60076 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_653
timestamp 1644511149
transform 1 0 61180 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_109_665
timestamp 1644511149
transform 1 0 62284 0 -1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_109_671
timestamp 1644511149
transform 1 0 62836 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_109_673
timestamp 1644511149
transform 1 0 63020 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_685
timestamp 1644511149
transform 1 0 64124 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_697
timestamp 1644511149
transform 1 0 65228 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_709
timestamp 1644511149
transform 1 0 66332 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_109_721
timestamp 1644511149
transform 1 0 67436 0 -1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_109_727
timestamp 1644511149
transform 1 0 67988 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_109_729
timestamp 1644511149
transform 1 0 68172 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_741
timestamp 1644511149
transform 1 0 69276 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_753
timestamp 1644511149
transform 1 0 70380 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_765
timestamp 1644511149
transform 1 0 71484 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_109_777
timestamp 1644511149
transform 1 0 72588 0 -1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_109_783
timestamp 1644511149
transform 1 0 73140 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_109_785
timestamp 1644511149
transform 1 0 73324 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_797
timestamp 1644511149
transform 1 0 74428 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_809
timestamp 1644511149
transform 1 0 75532 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_821
timestamp 1644511149
transform 1 0 76636 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_109_833
timestamp 1644511149
transform 1 0 77740 0 -1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_109_839
timestamp 1644511149
transform 1 0 78292 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_109_841
timestamp 1644511149
transform 1 0 78476 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_110_3
timestamp 1644511149
transform 1 0 1380 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_15
timestamp 1644511149
transform 1 0 2484 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_110_27
timestamp 1644511149
transform 1 0 3588 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_110_29
timestamp 1644511149
transform 1 0 3772 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_41
timestamp 1644511149
transform 1 0 4876 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_53
timestamp 1644511149
transform 1 0 5980 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_65
timestamp 1644511149
transform 1 0 7084 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_110_77
timestamp 1644511149
transform 1 0 8188 0 1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_110_83
timestamp 1644511149
transform 1 0 8740 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_110_85
timestamp 1644511149
transform 1 0 8924 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_97
timestamp 1644511149
transform 1 0 10028 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_109
timestamp 1644511149
transform 1 0 11132 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_121
timestamp 1644511149
transform 1 0 12236 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_110_133
timestamp 1644511149
transform 1 0 13340 0 1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_110_139
timestamp 1644511149
transform 1 0 13892 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_110_141
timestamp 1644511149
transform 1 0 14076 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_153
timestamp 1644511149
transform 1 0 15180 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_165
timestamp 1644511149
transform 1 0 16284 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_177
timestamp 1644511149
transform 1 0 17388 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_110_189
timestamp 1644511149
transform 1 0 18492 0 1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_110_195
timestamp 1644511149
transform 1 0 19044 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_110_197
timestamp 1644511149
transform 1 0 19228 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_209
timestamp 1644511149
transform 1 0 20332 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_221
timestamp 1644511149
transform 1 0 21436 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_233
timestamp 1644511149
transform 1 0 22540 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_110_245
timestamp 1644511149
transform 1 0 23644 0 1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_110_251
timestamp 1644511149
transform 1 0 24196 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_110_253
timestamp 1644511149
transform 1 0 24380 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_265
timestamp 1644511149
transform 1 0 25484 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_277
timestamp 1644511149
transform 1 0 26588 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_289
timestamp 1644511149
transform 1 0 27692 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_110_301
timestamp 1644511149
transform 1 0 28796 0 1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_110_307
timestamp 1644511149
transform 1 0 29348 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_110_309
timestamp 1644511149
transform 1 0 29532 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_321
timestamp 1644511149
transform 1 0 30636 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_333
timestamp 1644511149
transform 1 0 31740 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_345
timestamp 1644511149
transform 1 0 32844 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_110_357
timestamp 1644511149
transform 1 0 33948 0 1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_110_363
timestamp 1644511149
transform 1 0 34500 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_110_365
timestamp 1644511149
transform 1 0 34684 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_377
timestamp 1644511149
transform 1 0 35788 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_389
timestamp 1644511149
transform 1 0 36892 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_401
timestamp 1644511149
transform 1 0 37996 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_110_413
timestamp 1644511149
transform 1 0 39100 0 1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_110_419
timestamp 1644511149
transform 1 0 39652 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_110_421
timestamp 1644511149
transform 1 0 39836 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_433
timestamp 1644511149
transform 1 0 40940 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_445
timestamp 1644511149
transform 1 0 42044 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_457
timestamp 1644511149
transform 1 0 43148 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_110_469
timestamp 1644511149
transform 1 0 44252 0 1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_110_475
timestamp 1644511149
transform 1 0 44804 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_110_477
timestamp 1644511149
transform 1 0 44988 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_489
timestamp 1644511149
transform 1 0 46092 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_501
timestamp 1644511149
transform 1 0 47196 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_513
timestamp 1644511149
transform 1 0 48300 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_110_525
timestamp 1644511149
transform 1 0 49404 0 1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_110_531
timestamp 1644511149
transform 1 0 49956 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_110_533
timestamp 1644511149
transform 1 0 50140 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_545
timestamp 1644511149
transform 1 0 51244 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_557
timestamp 1644511149
transform 1 0 52348 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_569
timestamp 1644511149
transform 1 0 53452 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_110_581
timestamp 1644511149
transform 1 0 54556 0 1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_110_587
timestamp 1644511149
transform 1 0 55108 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_110_589
timestamp 1644511149
transform 1 0 55292 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_601
timestamp 1644511149
transform 1 0 56396 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_613
timestamp 1644511149
transform 1 0 57500 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_625
timestamp 1644511149
transform 1 0 58604 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_110_637
timestamp 1644511149
transform 1 0 59708 0 1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_110_643
timestamp 1644511149
transform 1 0 60260 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_110_645
timestamp 1644511149
transform 1 0 60444 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_657
timestamp 1644511149
transform 1 0 61548 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_669
timestamp 1644511149
transform 1 0 62652 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_681
timestamp 1644511149
transform 1 0 63756 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_110_693
timestamp 1644511149
transform 1 0 64860 0 1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_110_699
timestamp 1644511149
transform 1 0 65412 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_110_701
timestamp 1644511149
transform 1 0 65596 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_713
timestamp 1644511149
transform 1 0 66700 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_725
timestamp 1644511149
transform 1 0 67804 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_737
timestamp 1644511149
transform 1 0 68908 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_110_749
timestamp 1644511149
transform 1 0 70012 0 1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_110_755
timestamp 1644511149
transform 1 0 70564 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_110_757
timestamp 1644511149
transform 1 0 70748 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_769
timestamp 1644511149
transform 1 0 71852 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_781
timestamp 1644511149
transform 1 0 72956 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_793
timestamp 1644511149
transform 1 0 74060 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_110_805
timestamp 1644511149
transform 1 0 75164 0 1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_110_811
timestamp 1644511149
transform 1 0 75716 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_110_813
timestamp 1644511149
transform 1 0 75900 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_825
timestamp 1644511149
transform 1 0 77004 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_110_837
timestamp 1644511149
transform 1 0 78108 0 1 62016
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_110_841
timestamp 1644511149
transform 1 0 78476 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_111_7
timestamp 1644511149
transform 1 0 1748 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_19
timestamp 1644511149
transform 1 0 2852 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_31
timestamp 1644511149
transform 1 0 3956 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_43
timestamp 1644511149
transform 1 0 5060 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_111_55
timestamp 1644511149
transform 1 0 6164 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_111_57
timestamp 1644511149
transform 1 0 6348 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_69
timestamp 1644511149
transform 1 0 7452 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_81
timestamp 1644511149
transform 1 0 8556 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_93
timestamp 1644511149
transform 1 0 9660 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_111_105
timestamp 1644511149
transform 1 0 10764 0 -1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_111_111
timestamp 1644511149
transform 1 0 11316 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_111_113
timestamp 1644511149
transform 1 0 11500 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_125
timestamp 1644511149
transform 1 0 12604 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_137
timestamp 1644511149
transform 1 0 13708 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_149
timestamp 1644511149
transform 1 0 14812 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_111_161
timestamp 1644511149
transform 1 0 15916 0 -1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_111_167
timestamp 1644511149
transform 1 0 16468 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_111_169
timestamp 1644511149
transform 1 0 16652 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_181
timestamp 1644511149
transform 1 0 17756 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_193
timestamp 1644511149
transform 1 0 18860 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_205
timestamp 1644511149
transform 1 0 19964 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_111_217
timestamp 1644511149
transform 1 0 21068 0 -1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_111_223
timestamp 1644511149
transform 1 0 21620 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_111_225
timestamp 1644511149
transform 1 0 21804 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_237
timestamp 1644511149
transform 1 0 22908 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_249
timestamp 1644511149
transform 1 0 24012 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_261
timestamp 1644511149
transform 1 0 25116 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_111_273
timestamp 1644511149
transform 1 0 26220 0 -1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_111_279
timestamp 1644511149
transform 1 0 26772 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_111_281
timestamp 1644511149
transform 1 0 26956 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_293
timestamp 1644511149
transform 1 0 28060 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_305
timestamp 1644511149
transform 1 0 29164 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_317
timestamp 1644511149
transform 1 0 30268 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_111_329
timestamp 1644511149
transform 1 0 31372 0 -1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_111_335
timestamp 1644511149
transform 1 0 31924 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_111_337
timestamp 1644511149
transform 1 0 32108 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_349
timestamp 1644511149
transform 1 0 33212 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_361
timestamp 1644511149
transform 1 0 34316 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_373
timestamp 1644511149
transform 1 0 35420 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_111_385
timestamp 1644511149
transform 1 0 36524 0 -1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_111_391
timestamp 1644511149
transform 1 0 37076 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_111_393
timestamp 1644511149
transform 1 0 37260 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_405
timestamp 1644511149
transform 1 0 38364 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_417
timestamp 1644511149
transform 1 0 39468 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_429
timestamp 1644511149
transform 1 0 40572 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_111_441
timestamp 1644511149
transform 1 0 41676 0 -1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_111_447
timestamp 1644511149
transform 1 0 42228 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_111_449
timestamp 1644511149
transform 1 0 42412 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_461
timestamp 1644511149
transform 1 0 43516 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_473
timestamp 1644511149
transform 1 0 44620 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_485
timestamp 1644511149
transform 1 0 45724 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_111_497
timestamp 1644511149
transform 1 0 46828 0 -1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_111_503
timestamp 1644511149
transform 1 0 47380 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_111_505
timestamp 1644511149
transform 1 0 47564 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_517
timestamp 1644511149
transform 1 0 48668 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_529
timestamp 1644511149
transform 1 0 49772 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_541
timestamp 1644511149
transform 1 0 50876 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_111_553
timestamp 1644511149
transform 1 0 51980 0 -1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_111_559
timestamp 1644511149
transform 1 0 52532 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_111_561
timestamp 1644511149
transform 1 0 52716 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_573
timestamp 1644511149
transform 1 0 53820 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_585
timestamp 1644511149
transform 1 0 54924 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_597
timestamp 1644511149
transform 1 0 56028 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_111_609
timestamp 1644511149
transform 1 0 57132 0 -1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_111_615
timestamp 1644511149
transform 1 0 57684 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_111_617
timestamp 1644511149
transform 1 0 57868 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_629
timestamp 1644511149
transform 1 0 58972 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_641
timestamp 1644511149
transform 1 0 60076 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_653
timestamp 1644511149
transform 1 0 61180 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_111_665
timestamp 1644511149
transform 1 0 62284 0 -1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_111_671
timestamp 1644511149
transform 1 0 62836 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_111_673
timestamp 1644511149
transform 1 0 63020 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_685
timestamp 1644511149
transform 1 0 64124 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_697
timestamp 1644511149
transform 1 0 65228 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_709
timestamp 1644511149
transform 1 0 66332 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_111_721
timestamp 1644511149
transform 1 0 67436 0 -1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_111_727
timestamp 1644511149
transform 1 0 67988 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_111_729
timestamp 1644511149
transform 1 0 68172 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_741
timestamp 1644511149
transform 1 0 69276 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_753
timestamp 1644511149
transform 1 0 70380 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_765
timestamp 1644511149
transform 1 0 71484 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_111_777
timestamp 1644511149
transform 1 0 72588 0 -1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_111_783
timestamp 1644511149
transform 1 0 73140 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_111_785
timestamp 1644511149
transform 1 0 73324 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_797
timestamp 1644511149
transform 1 0 74428 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_809
timestamp 1644511149
transform 1 0 75532 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_821
timestamp 1644511149
transform 1 0 76636 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_111_833
timestamp 1644511149
transform 1 0 77740 0 -1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_111_839
timestamp 1644511149
transform 1 0 78292 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_111_841
timestamp 1644511149
transform 1 0 78476 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_112_3
timestamp 1644511149
transform 1 0 1380 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_15
timestamp 1644511149
transform 1 0 2484 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_112_27
timestamp 1644511149
transform 1 0 3588 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_112_29
timestamp 1644511149
transform 1 0 3772 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_41
timestamp 1644511149
transform 1 0 4876 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_53
timestamp 1644511149
transform 1 0 5980 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_65
timestamp 1644511149
transform 1 0 7084 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_112_77
timestamp 1644511149
transform 1 0 8188 0 1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_112_83
timestamp 1644511149
transform 1 0 8740 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_112_85
timestamp 1644511149
transform 1 0 8924 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_97
timestamp 1644511149
transform 1 0 10028 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_109
timestamp 1644511149
transform 1 0 11132 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_121
timestamp 1644511149
transform 1 0 12236 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_112_133
timestamp 1644511149
transform 1 0 13340 0 1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_112_139
timestamp 1644511149
transform 1 0 13892 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_112_141
timestamp 1644511149
transform 1 0 14076 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_153
timestamp 1644511149
transform 1 0 15180 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_165
timestamp 1644511149
transform 1 0 16284 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_177
timestamp 1644511149
transform 1 0 17388 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_112_189
timestamp 1644511149
transform 1 0 18492 0 1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_112_195
timestamp 1644511149
transform 1 0 19044 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_112_197
timestamp 1644511149
transform 1 0 19228 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_209
timestamp 1644511149
transform 1 0 20332 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_221
timestamp 1644511149
transform 1 0 21436 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_233
timestamp 1644511149
transform 1 0 22540 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_112_245
timestamp 1644511149
transform 1 0 23644 0 1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_112_251
timestamp 1644511149
transform 1 0 24196 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_112_253
timestamp 1644511149
transform 1 0 24380 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_265
timestamp 1644511149
transform 1 0 25484 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_277
timestamp 1644511149
transform 1 0 26588 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_289
timestamp 1644511149
transform 1 0 27692 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_112_301
timestamp 1644511149
transform 1 0 28796 0 1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_112_307
timestamp 1644511149
transform 1 0 29348 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_112_309
timestamp 1644511149
transform 1 0 29532 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_321
timestamp 1644511149
transform 1 0 30636 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_333
timestamp 1644511149
transform 1 0 31740 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_345
timestamp 1644511149
transform 1 0 32844 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_112_357
timestamp 1644511149
transform 1 0 33948 0 1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_112_363
timestamp 1644511149
transform 1 0 34500 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_112_365
timestamp 1644511149
transform 1 0 34684 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_377
timestamp 1644511149
transform 1 0 35788 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_389
timestamp 1644511149
transform 1 0 36892 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_401
timestamp 1644511149
transform 1 0 37996 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_112_413
timestamp 1644511149
transform 1 0 39100 0 1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_112_419
timestamp 1644511149
transform 1 0 39652 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_112_421
timestamp 1644511149
transform 1 0 39836 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_433
timestamp 1644511149
transform 1 0 40940 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_445
timestamp 1644511149
transform 1 0 42044 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_457
timestamp 1644511149
transform 1 0 43148 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_112_469
timestamp 1644511149
transform 1 0 44252 0 1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_112_475
timestamp 1644511149
transform 1 0 44804 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_112_477
timestamp 1644511149
transform 1 0 44988 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_489
timestamp 1644511149
transform 1 0 46092 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_501
timestamp 1644511149
transform 1 0 47196 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_513
timestamp 1644511149
transform 1 0 48300 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_112_525
timestamp 1644511149
transform 1 0 49404 0 1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_112_531
timestamp 1644511149
transform 1 0 49956 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_112_533
timestamp 1644511149
transform 1 0 50140 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_545
timestamp 1644511149
transform 1 0 51244 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_557
timestamp 1644511149
transform 1 0 52348 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_569
timestamp 1644511149
transform 1 0 53452 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_112_581
timestamp 1644511149
transform 1 0 54556 0 1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_112_587
timestamp 1644511149
transform 1 0 55108 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_112_589
timestamp 1644511149
transform 1 0 55292 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_601
timestamp 1644511149
transform 1 0 56396 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_613
timestamp 1644511149
transform 1 0 57500 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_625
timestamp 1644511149
transform 1 0 58604 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_112_637
timestamp 1644511149
transform 1 0 59708 0 1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_112_643
timestamp 1644511149
transform 1 0 60260 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_112_645
timestamp 1644511149
transform 1 0 60444 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_657
timestamp 1644511149
transform 1 0 61548 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_669
timestamp 1644511149
transform 1 0 62652 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_681
timestamp 1644511149
transform 1 0 63756 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_112_693
timestamp 1644511149
transform 1 0 64860 0 1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_112_699
timestamp 1644511149
transform 1 0 65412 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_112_701
timestamp 1644511149
transform 1 0 65596 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_713
timestamp 1644511149
transform 1 0 66700 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_725
timestamp 1644511149
transform 1 0 67804 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_737
timestamp 1644511149
transform 1 0 68908 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_112_749
timestamp 1644511149
transform 1 0 70012 0 1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_112_755
timestamp 1644511149
transform 1 0 70564 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_112_757
timestamp 1644511149
transform 1 0 70748 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_769
timestamp 1644511149
transform 1 0 71852 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_781
timestamp 1644511149
transform 1 0 72956 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_793
timestamp 1644511149
transform 1 0 74060 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_112_805
timestamp 1644511149
transform 1 0 75164 0 1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_112_811
timestamp 1644511149
transform 1 0 75716 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_112_813
timestamp 1644511149
transform 1 0 75900 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_112_825
timestamp 1644511149
transform 1 0 77004 0 1 63104
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_112_829
timestamp 1644511149
transform 1 0 77372 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_112_832
timestamp 1644511149
transform 1 0 77648 0 1 63104
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_112_838
timestamp 1644511149
transform 1 0 78200 0 1 63104
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_113_3
timestamp 1644511149
transform 1 0 1380 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_15
timestamp 1644511149
transform 1 0 2484 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_27
timestamp 1644511149
transform 1 0 3588 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_39
timestamp 1644511149
transform 1 0 4692 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_113_51
timestamp 1644511149
transform 1 0 5796 0 -1 64192
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_113_55
timestamp 1644511149
transform 1 0 6164 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_113_57
timestamp 1644511149
transform 1 0 6348 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_69
timestamp 1644511149
transform 1 0 7452 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_81
timestamp 1644511149
transform 1 0 8556 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_93
timestamp 1644511149
transform 1 0 9660 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_113_105
timestamp 1644511149
transform 1 0 10764 0 -1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_113_111
timestamp 1644511149
transform 1 0 11316 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_113_113
timestamp 1644511149
transform 1 0 11500 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_125
timestamp 1644511149
transform 1 0 12604 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_137
timestamp 1644511149
transform 1 0 13708 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_149
timestamp 1644511149
transform 1 0 14812 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_113_161
timestamp 1644511149
transform 1 0 15916 0 -1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_113_167
timestamp 1644511149
transform 1 0 16468 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_113_169
timestamp 1644511149
transform 1 0 16652 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_181
timestamp 1644511149
transform 1 0 17756 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_193
timestamp 1644511149
transform 1 0 18860 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_205
timestamp 1644511149
transform 1 0 19964 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_113_217
timestamp 1644511149
transform 1 0 21068 0 -1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_113_223
timestamp 1644511149
transform 1 0 21620 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_113_225
timestamp 1644511149
transform 1 0 21804 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_237
timestamp 1644511149
transform 1 0 22908 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_249
timestamp 1644511149
transform 1 0 24012 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_261
timestamp 1644511149
transform 1 0 25116 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_113_273
timestamp 1644511149
transform 1 0 26220 0 -1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_113_279
timestamp 1644511149
transform 1 0 26772 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_113_281
timestamp 1644511149
transform 1 0 26956 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_293
timestamp 1644511149
transform 1 0 28060 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_305
timestamp 1644511149
transform 1 0 29164 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_317
timestamp 1644511149
transform 1 0 30268 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_113_329
timestamp 1644511149
transform 1 0 31372 0 -1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_113_335
timestamp 1644511149
transform 1 0 31924 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_113_337
timestamp 1644511149
transform 1 0 32108 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_349
timestamp 1644511149
transform 1 0 33212 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_361
timestamp 1644511149
transform 1 0 34316 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_373
timestamp 1644511149
transform 1 0 35420 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_113_385
timestamp 1644511149
transform 1 0 36524 0 -1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_113_391
timestamp 1644511149
transform 1 0 37076 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_113_393
timestamp 1644511149
transform 1 0 37260 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_405
timestamp 1644511149
transform 1 0 38364 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_420
timestamp 1644511149
transform 1 0 39744 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_432
timestamp 1644511149
transform 1 0 40848 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_113_444
timestamp 1644511149
transform 1 0 41952 0 -1 64192
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_113_449
timestamp 1644511149
transform 1 0 42412 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_461
timestamp 1644511149
transform 1 0 43516 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_473
timestamp 1644511149
transform 1 0 44620 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_485
timestamp 1644511149
transform 1 0 45724 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_113_497
timestamp 1644511149
transform 1 0 46828 0 -1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_113_503
timestamp 1644511149
transform 1 0 47380 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_113_505
timestamp 1644511149
transform 1 0 47564 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_517
timestamp 1644511149
transform 1 0 48668 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_529
timestamp 1644511149
transform 1 0 49772 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_541
timestamp 1644511149
transform 1 0 50876 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_113_553
timestamp 1644511149
transform 1 0 51980 0 -1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_113_559
timestamp 1644511149
transform 1 0 52532 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_113_561
timestamp 1644511149
transform 1 0 52716 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_573
timestamp 1644511149
transform 1 0 53820 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_585
timestamp 1644511149
transform 1 0 54924 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_597
timestamp 1644511149
transform 1 0 56028 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_113_609
timestamp 1644511149
transform 1 0 57132 0 -1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_113_615
timestamp 1644511149
transform 1 0 57684 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_113_617
timestamp 1644511149
transform 1 0 57868 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_629
timestamp 1644511149
transform 1 0 58972 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_641
timestamp 1644511149
transform 1 0 60076 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_653
timestamp 1644511149
transform 1 0 61180 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_113_665
timestamp 1644511149
transform 1 0 62284 0 -1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_113_671
timestamp 1644511149
transform 1 0 62836 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_113_673
timestamp 1644511149
transform 1 0 63020 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_685
timestamp 1644511149
transform 1 0 64124 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_697
timestamp 1644511149
transform 1 0 65228 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_709
timestamp 1644511149
transform 1 0 66332 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_113_721
timestamp 1644511149
transform 1 0 67436 0 -1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_113_727
timestamp 1644511149
transform 1 0 67988 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_113_729
timestamp 1644511149
transform 1 0 68172 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_741
timestamp 1644511149
transform 1 0 69276 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_753
timestamp 1644511149
transform 1 0 70380 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_765
timestamp 1644511149
transform 1 0 71484 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_113_777
timestamp 1644511149
transform 1 0 72588 0 -1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_113_783
timestamp 1644511149
transform 1 0 73140 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_113_785
timestamp 1644511149
transform 1 0 73324 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_797
timestamp 1644511149
transform 1 0 74428 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_809
timestamp 1644511149
transform 1 0 75532 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_821
timestamp 1644511149
transform 1 0 76636 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_113_833
timestamp 1644511149
transform 1 0 77740 0 -1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_113_839
timestamp 1644511149
transform 1 0 78292 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_113_841
timestamp 1644511149
transform 1 0 78476 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_114_3
timestamp 1644511149
transform 1 0 1380 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_15
timestamp 1644511149
transform 1 0 2484 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_114_27
timestamp 1644511149
transform 1 0 3588 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_114_29
timestamp 1644511149
transform 1 0 3772 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_41
timestamp 1644511149
transform 1 0 4876 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_53
timestamp 1644511149
transform 1 0 5980 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_65
timestamp 1644511149
transform 1 0 7084 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_114_77
timestamp 1644511149
transform 1 0 8188 0 1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_114_83
timestamp 1644511149
transform 1 0 8740 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_114_85
timestamp 1644511149
transform 1 0 8924 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_97
timestamp 1644511149
transform 1 0 10028 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_109
timestamp 1644511149
transform 1 0 11132 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_121
timestamp 1644511149
transform 1 0 12236 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_114_133
timestamp 1644511149
transform 1 0 13340 0 1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_114_139
timestamp 1644511149
transform 1 0 13892 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_114_141
timestamp 1644511149
transform 1 0 14076 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_153
timestamp 1644511149
transform 1 0 15180 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_165
timestamp 1644511149
transform 1 0 16284 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_177
timestamp 1644511149
transform 1 0 17388 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_114_189
timestamp 1644511149
transform 1 0 18492 0 1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_114_195
timestamp 1644511149
transform 1 0 19044 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_114_197
timestamp 1644511149
transform 1 0 19228 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_209
timestamp 1644511149
transform 1 0 20332 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_221
timestamp 1644511149
transform 1 0 21436 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_233
timestamp 1644511149
transform 1 0 22540 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_114_245
timestamp 1644511149
transform 1 0 23644 0 1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_114_251
timestamp 1644511149
transform 1 0 24196 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_114_253
timestamp 1644511149
transform 1 0 24380 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_265
timestamp 1644511149
transform 1 0 25484 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_277
timestamp 1644511149
transform 1 0 26588 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_289
timestamp 1644511149
transform 1 0 27692 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_114_301
timestamp 1644511149
transform 1 0 28796 0 1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_114_307
timestamp 1644511149
transform 1 0 29348 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_114_309
timestamp 1644511149
transform 1 0 29532 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_321
timestamp 1644511149
transform 1 0 30636 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_333
timestamp 1644511149
transform 1 0 31740 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_345
timestamp 1644511149
transform 1 0 32844 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_114_357
timestamp 1644511149
transform 1 0 33948 0 1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_114_363
timestamp 1644511149
transform 1 0 34500 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_114_365
timestamp 1644511149
transform 1 0 34684 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_377
timestamp 1644511149
transform 1 0 35788 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_389
timestamp 1644511149
transform 1 0 36892 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_401
timestamp 1644511149
transform 1 0 37996 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_114_413
timestamp 1644511149
transform 1 0 39100 0 1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_114_419
timestamp 1644511149
transform 1 0 39652 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_114_421
timestamp 1644511149
transform 1 0 39836 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_114_438
timestamp 1644511149
transform 1 0 41400 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_450
timestamp 1644511149
transform 1 0 42504 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_462
timestamp 1644511149
transform 1 0 43608 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_114_474
timestamp 1644511149
transform 1 0 44712 0 1 64192
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_114_477
timestamp 1644511149
transform 1 0 44988 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_489
timestamp 1644511149
transform 1 0 46092 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_501
timestamp 1644511149
transform 1 0 47196 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_513
timestamp 1644511149
transform 1 0 48300 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_114_525
timestamp 1644511149
transform 1 0 49404 0 1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_114_531
timestamp 1644511149
transform 1 0 49956 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_114_533
timestamp 1644511149
transform 1 0 50140 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_545
timestamp 1644511149
transform 1 0 51244 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_557
timestamp 1644511149
transform 1 0 52348 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_569
timestamp 1644511149
transform 1 0 53452 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_114_581
timestamp 1644511149
transform 1 0 54556 0 1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_114_587
timestamp 1644511149
transform 1 0 55108 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_114_589
timestamp 1644511149
transform 1 0 55292 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_601
timestamp 1644511149
transform 1 0 56396 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_613
timestamp 1644511149
transform 1 0 57500 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_625
timestamp 1644511149
transform 1 0 58604 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_114_637
timestamp 1644511149
transform 1 0 59708 0 1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_114_643
timestamp 1644511149
transform 1 0 60260 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_114_645
timestamp 1644511149
transform 1 0 60444 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_657
timestamp 1644511149
transform 1 0 61548 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_669
timestamp 1644511149
transform 1 0 62652 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_681
timestamp 1644511149
transform 1 0 63756 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_114_693
timestamp 1644511149
transform 1 0 64860 0 1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_114_699
timestamp 1644511149
transform 1 0 65412 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_114_701
timestamp 1644511149
transform 1 0 65596 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_713
timestamp 1644511149
transform 1 0 66700 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_725
timestamp 1644511149
transform 1 0 67804 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_737
timestamp 1644511149
transform 1 0 68908 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_114_749
timestamp 1644511149
transform 1 0 70012 0 1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_114_755
timestamp 1644511149
transform 1 0 70564 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_114_757
timestamp 1644511149
transform 1 0 70748 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_769
timestamp 1644511149
transform 1 0 71852 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_781
timestamp 1644511149
transform 1 0 72956 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_793
timestamp 1644511149
transform 1 0 74060 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_114_805
timestamp 1644511149
transform 1 0 75164 0 1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_114_811
timestamp 1644511149
transform 1 0 75716 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_114_813
timestamp 1644511149
transform 1 0 75900 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_825
timestamp 1644511149
transform 1 0 77004 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_114_837
timestamp 1644511149
transform 1 0 78108 0 1 64192
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_114_841
timestamp 1644511149
transform 1 0 78476 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_115_3
timestamp 1644511149
transform 1 0 1380 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_15
timestamp 1644511149
transform 1 0 2484 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_27
timestamp 1644511149
transform 1 0 3588 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_39
timestamp 1644511149
transform 1 0 4692 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_115_51
timestamp 1644511149
transform 1 0 5796 0 -1 65280
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_115_55
timestamp 1644511149
transform 1 0 6164 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_115_57
timestamp 1644511149
transform 1 0 6348 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_69
timestamp 1644511149
transform 1 0 7452 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_81
timestamp 1644511149
transform 1 0 8556 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_93
timestamp 1644511149
transform 1 0 9660 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_115_105
timestamp 1644511149
transform 1 0 10764 0 -1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_115_111
timestamp 1644511149
transform 1 0 11316 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_115_113
timestamp 1644511149
transform 1 0 11500 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_125
timestamp 1644511149
transform 1 0 12604 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_137
timestamp 1644511149
transform 1 0 13708 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_149
timestamp 1644511149
transform 1 0 14812 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_115_161
timestamp 1644511149
transform 1 0 15916 0 -1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_115_167
timestamp 1644511149
transform 1 0 16468 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_115_169
timestamp 1644511149
transform 1 0 16652 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_181
timestamp 1644511149
transform 1 0 17756 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_193
timestamp 1644511149
transform 1 0 18860 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_205
timestamp 1644511149
transform 1 0 19964 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_115_217
timestamp 1644511149
transform 1 0 21068 0 -1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_115_223
timestamp 1644511149
transform 1 0 21620 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_115_225
timestamp 1644511149
transform 1 0 21804 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_237
timestamp 1644511149
transform 1 0 22908 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_249
timestamp 1644511149
transform 1 0 24012 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_261
timestamp 1644511149
transform 1 0 25116 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_115_273
timestamp 1644511149
transform 1 0 26220 0 -1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_115_279
timestamp 1644511149
transform 1 0 26772 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_115_281
timestamp 1644511149
transform 1 0 26956 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_293
timestamp 1644511149
transform 1 0 28060 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_305
timestamp 1644511149
transform 1 0 29164 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_317
timestamp 1644511149
transform 1 0 30268 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_115_329
timestamp 1644511149
transform 1 0 31372 0 -1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_115_335
timestamp 1644511149
transform 1 0 31924 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_115_337
timestamp 1644511149
transform 1 0 32108 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_349
timestamp 1644511149
transform 1 0 33212 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_361
timestamp 1644511149
transform 1 0 34316 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_373
timestamp 1644511149
transform 1 0 35420 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_115_385
timestamp 1644511149
transform 1 0 36524 0 -1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_115_391
timestamp 1644511149
transform 1 0 37076 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_115_393
timestamp 1644511149
transform 1 0 37260 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_405
timestamp 1644511149
transform 1 0 38364 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_115_417
timestamp 1644511149
transform 1 0 39468 0 -1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_115_426
timestamp 1644511149
transform 1 0 40296 0 -1 65280
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_115_437
timestamp 1644511149
transform 1 0 41308 0 -1 65280
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_115_445
timestamp 1644511149
transform 1 0 42044 0 -1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_115_449
timestamp 1644511149
transform 1 0 42412 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_461
timestamp 1644511149
transform 1 0 43516 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_473
timestamp 1644511149
transform 1 0 44620 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_485
timestamp 1644511149
transform 1 0 45724 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_115_497
timestamp 1644511149
transform 1 0 46828 0 -1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_115_503
timestamp 1644511149
transform 1 0 47380 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_115_505
timestamp 1644511149
transform 1 0 47564 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_517
timestamp 1644511149
transform 1 0 48668 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_529
timestamp 1644511149
transform 1 0 49772 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_541
timestamp 1644511149
transform 1 0 50876 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_115_553
timestamp 1644511149
transform 1 0 51980 0 -1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_115_559
timestamp 1644511149
transform 1 0 52532 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_115_561
timestamp 1644511149
transform 1 0 52716 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_573
timestamp 1644511149
transform 1 0 53820 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_585
timestamp 1644511149
transform 1 0 54924 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_597
timestamp 1644511149
transform 1 0 56028 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_115_609
timestamp 1644511149
transform 1 0 57132 0 -1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_115_615
timestamp 1644511149
transform 1 0 57684 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_115_617
timestamp 1644511149
transform 1 0 57868 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_629
timestamp 1644511149
transform 1 0 58972 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_641
timestamp 1644511149
transform 1 0 60076 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_653
timestamp 1644511149
transform 1 0 61180 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_115_665
timestamp 1644511149
transform 1 0 62284 0 -1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_115_671
timestamp 1644511149
transform 1 0 62836 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_115_673
timestamp 1644511149
transform 1 0 63020 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_685
timestamp 1644511149
transform 1 0 64124 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_697
timestamp 1644511149
transform 1 0 65228 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_709
timestamp 1644511149
transform 1 0 66332 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_115_721
timestamp 1644511149
transform 1 0 67436 0 -1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_115_727
timestamp 1644511149
transform 1 0 67988 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_115_729
timestamp 1644511149
transform 1 0 68172 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_741
timestamp 1644511149
transform 1 0 69276 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_753
timestamp 1644511149
transform 1 0 70380 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_765
timestamp 1644511149
transform 1 0 71484 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_115_777
timestamp 1644511149
transform 1 0 72588 0 -1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_115_783
timestamp 1644511149
transform 1 0 73140 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_115_785
timestamp 1644511149
transform 1 0 73324 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_797
timestamp 1644511149
transform 1 0 74428 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_809
timestamp 1644511149
transform 1 0 75532 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_821
timestamp 1644511149
transform 1 0 76636 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_115_833
timestamp 1644511149
transform 1 0 77740 0 -1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_115_839
timestamp 1644511149
transform 1 0 78292 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_115_841
timestamp 1644511149
transform 1 0 78476 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_116_3
timestamp 1644511149
transform 1 0 1380 0 1 65280
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_116_11
timestamp 1644511149
transform 1 0 2116 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_116_23
timestamp 1644511149
transform 1 0 3220 0 1 65280
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_116_27
timestamp 1644511149
transform 1 0 3588 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_116_29
timestamp 1644511149
transform 1 0 3772 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_41
timestamp 1644511149
transform 1 0 4876 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_53
timestamp 1644511149
transform 1 0 5980 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_65
timestamp 1644511149
transform 1 0 7084 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_116_77
timestamp 1644511149
transform 1 0 8188 0 1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_116_83
timestamp 1644511149
transform 1 0 8740 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_116_85
timestamp 1644511149
transform 1 0 8924 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_97
timestamp 1644511149
transform 1 0 10028 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_109
timestamp 1644511149
transform 1 0 11132 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_121
timestamp 1644511149
transform 1 0 12236 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_116_133
timestamp 1644511149
transform 1 0 13340 0 1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_116_139
timestamp 1644511149
transform 1 0 13892 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_116_141
timestamp 1644511149
transform 1 0 14076 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_153
timestamp 1644511149
transform 1 0 15180 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_165
timestamp 1644511149
transform 1 0 16284 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_177
timestamp 1644511149
transform 1 0 17388 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_116_189
timestamp 1644511149
transform 1 0 18492 0 1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_116_195
timestamp 1644511149
transform 1 0 19044 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_116_197
timestamp 1644511149
transform 1 0 19228 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_209
timestamp 1644511149
transform 1 0 20332 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_221
timestamp 1644511149
transform 1 0 21436 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_233
timestamp 1644511149
transform 1 0 22540 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_116_245
timestamp 1644511149
transform 1 0 23644 0 1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_116_251
timestamp 1644511149
transform 1 0 24196 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_116_253
timestamp 1644511149
transform 1 0 24380 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_265
timestamp 1644511149
transform 1 0 25484 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_277
timestamp 1644511149
transform 1 0 26588 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_289
timestamp 1644511149
transform 1 0 27692 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_116_301
timestamp 1644511149
transform 1 0 28796 0 1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_116_307
timestamp 1644511149
transform 1 0 29348 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_116_309
timestamp 1644511149
transform 1 0 29532 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_321
timestamp 1644511149
transform 1 0 30636 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_333
timestamp 1644511149
transform 1 0 31740 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_345
timestamp 1644511149
transform 1 0 32844 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_116_357
timestamp 1644511149
transform 1 0 33948 0 1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_116_363
timestamp 1644511149
transform 1 0 34500 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_116_365
timestamp 1644511149
transform 1 0 34684 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_377
timestamp 1644511149
transform 1 0 35788 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_389
timestamp 1644511149
transform 1 0 36892 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_401
timestamp 1644511149
transform 1 0 37996 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_116_413
timestamp 1644511149
transform 1 0 39100 0 1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_116_419
timestamp 1644511149
transform 1 0 39652 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_116_444
timestamp 1644511149
transform 1 0 41952 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_456
timestamp 1644511149
transform 1 0 43056 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_116_468
timestamp 1644511149
transform 1 0 44160 0 1 65280
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_116_477
timestamp 1644511149
transform 1 0 44988 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_489
timestamp 1644511149
transform 1 0 46092 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_501
timestamp 1644511149
transform 1 0 47196 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_513
timestamp 1644511149
transform 1 0 48300 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_116_525
timestamp 1644511149
transform 1 0 49404 0 1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_116_531
timestamp 1644511149
transform 1 0 49956 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_116_533
timestamp 1644511149
transform 1 0 50140 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_545
timestamp 1644511149
transform 1 0 51244 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_557
timestamp 1644511149
transform 1 0 52348 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_569
timestamp 1644511149
transform 1 0 53452 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_116_581
timestamp 1644511149
transform 1 0 54556 0 1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_116_587
timestamp 1644511149
transform 1 0 55108 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_116_589
timestamp 1644511149
transform 1 0 55292 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_601
timestamp 1644511149
transform 1 0 56396 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_613
timestamp 1644511149
transform 1 0 57500 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_625
timestamp 1644511149
transform 1 0 58604 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_116_637
timestamp 1644511149
transform 1 0 59708 0 1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_116_643
timestamp 1644511149
transform 1 0 60260 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_116_645
timestamp 1644511149
transform 1 0 60444 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_657
timestamp 1644511149
transform 1 0 61548 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_669
timestamp 1644511149
transform 1 0 62652 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_681
timestamp 1644511149
transform 1 0 63756 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_116_693
timestamp 1644511149
transform 1 0 64860 0 1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_116_699
timestamp 1644511149
transform 1 0 65412 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_116_701
timestamp 1644511149
transform 1 0 65596 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_713
timestamp 1644511149
transform 1 0 66700 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_725
timestamp 1644511149
transform 1 0 67804 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_737
timestamp 1644511149
transform 1 0 68908 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_116_749
timestamp 1644511149
transform 1 0 70012 0 1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_116_755
timestamp 1644511149
transform 1 0 70564 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_116_757
timestamp 1644511149
transform 1 0 70748 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_769
timestamp 1644511149
transform 1 0 71852 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_781
timestamp 1644511149
transform 1 0 72956 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_793
timestamp 1644511149
transform 1 0 74060 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_116_805
timestamp 1644511149
transform 1 0 75164 0 1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_116_811
timestamp 1644511149
transform 1 0 75716 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_116_813
timestamp 1644511149
transform 1 0 75900 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_825
timestamp 1644511149
transform 1 0 77004 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_116_837
timestamp 1644511149
transform 1 0 78108 0 1 65280
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_116_841
timestamp 1644511149
transform 1 0 78476 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_117_7
timestamp 1644511149
transform 1 0 1748 0 -1 66368
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_117_14
timestamp 1644511149
transform 1 0 2392 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_26
timestamp 1644511149
transform 1 0 3496 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_38
timestamp 1644511149
transform 1 0 4600 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_117_50
timestamp 1644511149
transform 1 0 5704 0 -1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_117_57
timestamp 1644511149
transform 1 0 6348 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_69
timestamp 1644511149
transform 1 0 7452 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_81
timestamp 1644511149
transform 1 0 8556 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_93
timestamp 1644511149
transform 1 0 9660 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_117_105
timestamp 1644511149
transform 1 0 10764 0 -1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_117_111
timestamp 1644511149
transform 1 0 11316 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_117_113
timestamp 1644511149
transform 1 0 11500 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_125
timestamp 1644511149
transform 1 0 12604 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_137
timestamp 1644511149
transform 1 0 13708 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_149
timestamp 1644511149
transform 1 0 14812 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_117_161
timestamp 1644511149
transform 1 0 15916 0 -1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_117_167
timestamp 1644511149
transform 1 0 16468 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_117_169
timestamp 1644511149
transform 1 0 16652 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_181
timestamp 1644511149
transform 1 0 17756 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_193
timestamp 1644511149
transform 1 0 18860 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_205
timestamp 1644511149
transform 1 0 19964 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_117_217
timestamp 1644511149
transform 1 0 21068 0 -1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_117_223
timestamp 1644511149
transform 1 0 21620 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_117_225
timestamp 1644511149
transform 1 0 21804 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_237
timestamp 1644511149
transform 1 0 22908 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_249
timestamp 1644511149
transform 1 0 24012 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_261
timestamp 1644511149
transform 1 0 25116 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_117_273
timestamp 1644511149
transform 1 0 26220 0 -1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_117_279
timestamp 1644511149
transform 1 0 26772 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_117_281
timestamp 1644511149
transform 1 0 26956 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_293
timestamp 1644511149
transform 1 0 28060 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_305
timestamp 1644511149
transform 1 0 29164 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_317
timestamp 1644511149
transform 1 0 30268 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_117_329
timestamp 1644511149
transform 1 0 31372 0 -1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_117_335
timestamp 1644511149
transform 1 0 31924 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_117_337
timestamp 1644511149
transform 1 0 32108 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_349
timestamp 1644511149
transform 1 0 33212 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_361
timestamp 1644511149
transform 1 0 34316 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_373
timestamp 1644511149
transform 1 0 35420 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_117_385
timestamp 1644511149
transform 1 0 36524 0 -1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_117_391
timestamp 1644511149
transform 1 0 37076 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_117_393
timestamp 1644511149
transform 1 0 37260 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_405
timestamp 1644511149
transform 1 0 38364 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_417
timestamp 1644511149
transform 1 0 39468 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_429
timestamp 1644511149
transform 1 0 40572 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_117_441
timestamp 1644511149
transform 1 0 41676 0 -1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_117_447
timestamp 1644511149
transform 1 0 42228 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_117_449
timestamp 1644511149
transform 1 0 42412 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_461
timestamp 1644511149
transform 1 0 43516 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_473
timestamp 1644511149
transform 1 0 44620 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_485
timestamp 1644511149
transform 1 0 45724 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_117_497
timestamp 1644511149
transform 1 0 46828 0 -1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_117_503
timestamp 1644511149
transform 1 0 47380 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_117_505
timestamp 1644511149
transform 1 0 47564 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_517
timestamp 1644511149
transform 1 0 48668 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_529
timestamp 1644511149
transform 1 0 49772 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_541
timestamp 1644511149
transform 1 0 50876 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_117_553
timestamp 1644511149
transform 1 0 51980 0 -1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_117_559
timestamp 1644511149
transform 1 0 52532 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_117_561
timestamp 1644511149
transform 1 0 52716 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_573
timestamp 1644511149
transform 1 0 53820 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_585
timestamp 1644511149
transform 1 0 54924 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_597
timestamp 1644511149
transform 1 0 56028 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_117_609
timestamp 1644511149
transform 1 0 57132 0 -1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_117_615
timestamp 1644511149
transform 1 0 57684 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_117_617
timestamp 1644511149
transform 1 0 57868 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_629
timestamp 1644511149
transform 1 0 58972 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_641
timestamp 1644511149
transform 1 0 60076 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_653
timestamp 1644511149
transform 1 0 61180 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_117_665
timestamp 1644511149
transform 1 0 62284 0 -1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_117_671
timestamp 1644511149
transform 1 0 62836 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_117_673
timestamp 1644511149
transform 1 0 63020 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_685
timestamp 1644511149
transform 1 0 64124 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_697
timestamp 1644511149
transform 1 0 65228 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_709
timestamp 1644511149
transform 1 0 66332 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_117_721
timestamp 1644511149
transform 1 0 67436 0 -1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_117_727
timestamp 1644511149
transform 1 0 67988 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_117_729
timestamp 1644511149
transform 1 0 68172 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_741
timestamp 1644511149
transform 1 0 69276 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_753
timestamp 1644511149
transform 1 0 70380 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_765
timestamp 1644511149
transform 1 0 71484 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_117_777
timestamp 1644511149
transform 1 0 72588 0 -1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_117_783
timestamp 1644511149
transform 1 0 73140 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_117_785
timestamp 1644511149
transform 1 0 73324 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_797
timestamp 1644511149
transform 1 0 74428 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_809
timestamp 1644511149
transform 1 0 75532 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_821
timestamp 1644511149
transform 1 0 76636 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_117_833
timestamp 1644511149
transform 1 0 77740 0 -1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_117_839
timestamp 1644511149
transform 1 0 78292 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_117_841
timestamp 1644511149
transform 1 0 78476 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_118_3
timestamp 1644511149
transform 1 0 1380 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_15
timestamp 1644511149
transform 1 0 2484 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_118_27
timestamp 1644511149
transform 1 0 3588 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_118_29
timestamp 1644511149
transform 1 0 3772 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_41
timestamp 1644511149
transform 1 0 4876 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_53
timestamp 1644511149
transform 1 0 5980 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_65
timestamp 1644511149
transform 1 0 7084 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_77
timestamp 1644511149
transform 1 0 8188 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_118_83
timestamp 1644511149
transform 1 0 8740 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_118_85
timestamp 1644511149
transform 1 0 8924 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_97
timestamp 1644511149
transform 1 0 10028 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_109
timestamp 1644511149
transform 1 0 11132 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_121
timestamp 1644511149
transform 1 0 12236 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_133
timestamp 1644511149
transform 1 0 13340 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_118_139
timestamp 1644511149
transform 1 0 13892 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_118_141
timestamp 1644511149
transform 1 0 14076 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_153
timestamp 1644511149
transform 1 0 15180 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_165
timestamp 1644511149
transform 1 0 16284 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_177
timestamp 1644511149
transform 1 0 17388 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_189
timestamp 1644511149
transform 1 0 18492 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_118_195
timestamp 1644511149
transform 1 0 19044 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_118_197
timestamp 1644511149
transform 1 0 19228 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_209
timestamp 1644511149
transform 1 0 20332 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_221
timestamp 1644511149
transform 1 0 21436 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_233
timestamp 1644511149
transform 1 0 22540 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_245
timestamp 1644511149
transform 1 0 23644 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_118_251
timestamp 1644511149
transform 1 0 24196 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_118_253
timestamp 1644511149
transform 1 0 24380 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_265
timestamp 1644511149
transform 1 0 25484 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_277
timestamp 1644511149
transform 1 0 26588 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_289
timestamp 1644511149
transform 1 0 27692 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_301
timestamp 1644511149
transform 1 0 28796 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_118_307
timestamp 1644511149
transform 1 0 29348 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_118_309
timestamp 1644511149
transform 1 0 29532 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_321
timestamp 1644511149
transform 1 0 30636 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_333
timestamp 1644511149
transform 1 0 31740 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_345
timestamp 1644511149
transform 1 0 32844 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_357
timestamp 1644511149
transform 1 0 33948 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_118_363
timestamp 1644511149
transform 1 0 34500 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_118_365
timestamp 1644511149
transform 1 0 34684 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_377
timestamp 1644511149
transform 1 0 35788 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_389
timestamp 1644511149
transform 1 0 36892 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_401
timestamp 1644511149
transform 1 0 37996 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_413
timestamp 1644511149
transform 1 0 39100 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_118_419
timestamp 1644511149
transform 1 0 39652 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_118_421
timestamp 1644511149
transform 1 0 39836 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_433
timestamp 1644511149
transform 1 0 40940 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_445
timestamp 1644511149
transform 1 0 42044 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_457
timestamp 1644511149
transform 1 0 43148 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_469
timestamp 1644511149
transform 1 0 44252 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_118_475
timestamp 1644511149
transform 1 0 44804 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_118_477
timestamp 1644511149
transform 1 0 44988 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_489
timestamp 1644511149
transform 1 0 46092 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_501
timestamp 1644511149
transform 1 0 47196 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_513
timestamp 1644511149
transform 1 0 48300 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_525
timestamp 1644511149
transform 1 0 49404 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_118_531
timestamp 1644511149
transform 1 0 49956 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_118_533
timestamp 1644511149
transform 1 0 50140 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_545
timestamp 1644511149
transform 1 0 51244 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_557
timestamp 1644511149
transform 1 0 52348 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_569
timestamp 1644511149
transform 1 0 53452 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_581
timestamp 1644511149
transform 1 0 54556 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_118_587
timestamp 1644511149
transform 1 0 55108 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_118_589
timestamp 1644511149
transform 1 0 55292 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_601
timestamp 1644511149
transform 1 0 56396 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_613
timestamp 1644511149
transform 1 0 57500 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_625
timestamp 1644511149
transform 1 0 58604 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_637
timestamp 1644511149
transform 1 0 59708 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_118_643
timestamp 1644511149
transform 1 0 60260 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_118_645
timestamp 1644511149
transform 1 0 60444 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_657
timestamp 1644511149
transform 1 0 61548 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_669
timestamp 1644511149
transform 1 0 62652 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_681
timestamp 1644511149
transform 1 0 63756 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_693
timestamp 1644511149
transform 1 0 64860 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_118_699
timestamp 1644511149
transform 1 0 65412 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_118_701
timestamp 1644511149
transform 1 0 65596 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_713
timestamp 1644511149
transform 1 0 66700 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_725
timestamp 1644511149
transform 1 0 67804 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_737
timestamp 1644511149
transform 1 0 68908 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_749
timestamp 1644511149
transform 1 0 70012 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_118_755
timestamp 1644511149
transform 1 0 70564 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_118_757
timestamp 1644511149
transform 1 0 70748 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_769
timestamp 1644511149
transform 1 0 71852 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_781
timestamp 1644511149
transform 1 0 72956 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_793
timestamp 1644511149
transform 1 0 74060 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_805
timestamp 1644511149
transform 1 0 75164 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_118_811
timestamp 1644511149
transform 1 0 75716 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_118_813
timestamp 1644511149
transform 1 0 75900 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_825
timestamp 1644511149
transform 1 0 77004 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_118_837
timestamp 1644511149
transform 1 0 78108 0 1 66368
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_118_841
timestamp 1644511149
transform 1 0 78476 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_119_3
timestamp 1644511149
transform 1 0 1380 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_15
timestamp 1644511149
transform 1 0 2484 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_27
timestamp 1644511149
transform 1 0 3588 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_39
timestamp 1644511149
transform 1 0 4692 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_119_51
timestamp 1644511149
transform 1 0 5796 0 -1 67456
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_119_55
timestamp 1644511149
transform 1 0 6164 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_119_57
timestamp 1644511149
transform 1 0 6348 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_69
timestamp 1644511149
transform 1 0 7452 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_81
timestamp 1644511149
transform 1 0 8556 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_93
timestamp 1644511149
transform 1 0 9660 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_119_105
timestamp 1644511149
transform 1 0 10764 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_119_111
timestamp 1644511149
transform 1 0 11316 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_119_113
timestamp 1644511149
transform 1 0 11500 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_125
timestamp 1644511149
transform 1 0 12604 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_137
timestamp 1644511149
transform 1 0 13708 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_149
timestamp 1644511149
transform 1 0 14812 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_119_161
timestamp 1644511149
transform 1 0 15916 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_119_167
timestamp 1644511149
transform 1 0 16468 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_119_169
timestamp 1644511149
transform 1 0 16652 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_181
timestamp 1644511149
transform 1 0 17756 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_193
timestamp 1644511149
transform 1 0 18860 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_205
timestamp 1644511149
transform 1 0 19964 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_119_217
timestamp 1644511149
transform 1 0 21068 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_119_223
timestamp 1644511149
transform 1 0 21620 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_119_225
timestamp 1644511149
transform 1 0 21804 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_237
timestamp 1644511149
transform 1 0 22908 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_249
timestamp 1644511149
transform 1 0 24012 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_261
timestamp 1644511149
transform 1 0 25116 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_119_273
timestamp 1644511149
transform 1 0 26220 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_119_279
timestamp 1644511149
transform 1 0 26772 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_119_281
timestamp 1644511149
transform 1 0 26956 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_293
timestamp 1644511149
transform 1 0 28060 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_305
timestamp 1644511149
transform 1 0 29164 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_317
timestamp 1644511149
transform 1 0 30268 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_119_329
timestamp 1644511149
transform 1 0 31372 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_119_335
timestamp 1644511149
transform 1 0 31924 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_119_337
timestamp 1644511149
transform 1 0 32108 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_349
timestamp 1644511149
transform 1 0 33212 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_361
timestamp 1644511149
transform 1 0 34316 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_373
timestamp 1644511149
transform 1 0 35420 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_119_385
timestamp 1644511149
transform 1 0 36524 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_119_391
timestamp 1644511149
transform 1 0 37076 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_119_393
timestamp 1644511149
transform 1 0 37260 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_405
timestamp 1644511149
transform 1 0 38364 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_417
timestamp 1644511149
transform 1 0 39468 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_429
timestamp 1644511149
transform 1 0 40572 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_119_441
timestamp 1644511149
transform 1 0 41676 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_119_447
timestamp 1644511149
transform 1 0 42228 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_119_449
timestamp 1644511149
transform 1 0 42412 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_461
timestamp 1644511149
transform 1 0 43516 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_473
timestamp 1644511149
transform 1 0 44620 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_485
timestamp 1644511149
transform 1 0 45724 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_119_497
timestamp 1644511149
transform 1 0 46828 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_119_503
timestamp 1644511149
transform 1 0 47380 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_119_505
timestamp 1644511149
transform 1 0 47564 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_517
timestamp 1644511149
transform 1 0 48668 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_529
timestamp 1644511149
transform 1 0 49772 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_541
timestamp 1644511149
transform 1 0 50876 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_119_553
timestamp 1644511149
transform 1 0 51980 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_119_559
timestamp 1644511149
transform 1 0 52532 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_119_561
timestamp 1644511149
transform 1 0 52716 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_573
timestamp 1644511149
transform 1 0 53820 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_585
timestamp 1644511149
transform 1 0 54924 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_597
timestamp 1644511149
transform 1 0 56028 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_119_609
timestamp 1644511149
transform 1 0 57132 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_119_615
timestamp 1644511149
transform 1 0 57684 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_119_617
timestamp 1644511149
transform 1 0 57868 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_629
timestamp 1644511149
transform 1 0 58972 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_641
timestamp 1644511149
transform 1 0 60076 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_653
timestamp 1644511149
transform 1 0 61180 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_119_665
timestamp 1644511149
transform 1 0 62284 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_119_671
timestamp 1644511149
transform 1 0 62836 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_119_673
timestamp 1644511149
transform 1 0 63020 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_685
timestamp 1644511149
transform 1 0 64124 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_697
timestamp 1644511149
transform 1 0 65228 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_709
timestamp 1644511149
transform 1 0 66332 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_119_721
timestamp 1644511149
transform 1 0 67436 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_119_727
timestamp 1644511149
transform 1 0 67988 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_119_729
timestamp 1644511149
transform 1 0 68172 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_741
timestamp 1644511149
transform 1 0 69276 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_753
timestamp 1644511149
transform 1 0 70380 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_765
timestamp 1644511149
transform 1 0 71484 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_119_777
timestamp 1644511149
transform 1 0 72588 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_119_783
timestamp 1644511149
transform 1 0 73140 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_119_785
timestamp 1644511149
transform 1 0 73324 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_797
timestamp 1644511149
transform 1 0 74428 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_809
timestamp 1644511149
transform 1 0 75532 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_821
timestamp 1644511149
transform 1 0 76636 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_119_833
timestamp 1644511149
transform 1 0 77740 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_119_839
timestamp 1644511149
transform 1 0 78292 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_119_841
timestamp 1644511149
transform 1 0 78476 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_120_3
timestamp 1644511149
transform 1 0 1380 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_15
timestamp 1644511149
transform 1 0 2484 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_120_27
timestamp 1644511149
transform 1 0 3588 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_120_29
timestamp 1644511149
transform 1 0 3772 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_41
timestamp 1644511149
transform 1 0 4876 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_53
timestamp 1644511149
transform 1 0 5980 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_65
timestamp 1644511149
transform 1 0 7084 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_120_77
timestamp 1644511149
transform 1 0 8188 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_120_83
timestamp 1644511149
transform 1 0 8740 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_120_85
timestamp 1644511149
transform 1 0 8924 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_97
timestamp 1644511149
transform 1 0 10028 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_109
timestamp 1644511149
transform 1 0 11132 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_121
timestamp 1644511149
transform 1 0 12236 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_120_133
timestamp 1644511149
transform 1 0 13340 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_120_139
timestamp 1644511149
transform 1 0 13892 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_120_141
timestamp 1644511149
transform 1 0 14076 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_153
timestamp 1644511149
transform 1 0 15180 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_165
timestamp 1644511149
transform 1 0 16284 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_177
timestamp 1644511149
transform 1 0 17388 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_120_189
timestamp 1644511149
transform 1 0 18492 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_120_195
timestamp 1644511149
transform 1 0 19044 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_120_197
timestamp 1644511149
transform 1 0 19228 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_209
timestamp 1644511149
transform 1 0 20332 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_221
timestamp 1644511149
transform 1 0 21436 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_233
timestamp 1644511149
transform 1 0 22540 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_120_245
timestamp 1644511149
transform 1 0 23644 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_120_251
timestamp 1644511149
transform 1 0 24196 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_120_253
timestamp 1644511149
transform 1 0 24380 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_265
timestamp 1644511149
transform 1 0 25484 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_277
timestamp 1644511149
transform 1 0 26588 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_289
timestamp 1644511149
transform 1 0 27692 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_120_301
timestamp 1644511149
transform 1 0 28796 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_120_307
timestamp 1644511149
transform 1 0 29348 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_120_309
timestamp 1644511149
transform 1 0 29532 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_321
timestamp 1644511149
transform 1 0 30636 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_333
timestamp 1644511149
transform 1 0 31740 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_345
timestamp 1644511149
transform 1 0 32844 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_120_357
timestamp 1644511149
transform 1 0 33948 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_120_363
timestamp 1644511149
transform 1 0 34500 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_120_365
timestamp 1644511149
transform 1 0 34684 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_377
timestamp 1644511149
transform 1 0 35788 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_389
timestamp 1644511149
transform 1 0 36892 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_401
timestamp 1644511149
transform 1 0 37996 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_120_413
timestamp 1644511149
transform 1 0 39100 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_120_419
timestamp 1644511149
transform 1 0 39652 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_120_421
timestamp 1644511149
transform 1 0 39836 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_433
timestamp 1644511149
transform 1 0 40940 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_445
timestamp 1644511149
transform 1 0 42044 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_457
timestamp 1644511149
transform 1 0 43148 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_120_469
timestamp 1644511149
transform 1 0 44252 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_120_475
timestamp 1644511149
transform 1 0 44804 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_120_477
timestamp 1644511149
transform 1 0 44988 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_489
timestamp 1644511149
transform 1 0 46092 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_501
timestamp 1644511149
transform 1 0 47196 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_513
timestamp 1644511149
transform 1 0 48300 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_120_525
timestamp 1644511149
transform 1 0 49404 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_120_531
timestamp 1644511149
transform 1 0 49956 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_120_533
timestamp 1644511149
transform 1 0 50140 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_545
timestamp 1644511149
transform 1 0 51244 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_557
timestamp 1644511149
transform 1 0 52348 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_569
timestamp 1644511149
transform 1 0 53452 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_120_581
timestamp 1644511149
transform 1 0 54556 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_120_587
timestamp 1644511149
transform 1 0 55108 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_120_589
timestamp 1644511149
transform 1 0 55292 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_601
timestamp 1644511149
transform 1 0 56396 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_613
timestamp 1644511149
transform 1 0 57500 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_625
timestamp 1644511149
transform 1 0 58604 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_120_637
timestamp 1644511149
transform 1 0 59708 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_120_643
timestamp 1644511149
transform 1 0 60260 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_120_645
timestamp 1644511149
transform 1 0 60444 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_657
timestamp 1644511149
transform 1 0 61548 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_669
timestamp 1644511149
transform 1 0 62652 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_681
timestamp 1644511149
transform 1 0 63756 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_120_693
timestamp 1644511149
transform 1 0 64860 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_120_699
timestamp 1644511149
transform 1 0 65412 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_120_701
timestamp 1644511149
transform 1 0 65596 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_713
timestamp 1644511149
transform 1 0 66700 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_725
timestamp 1644511149
transform 1 0 67804 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_737
timestamp 1644511149
transform 1 0 68908 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_120_749
timestamp 1644511149
transform 1 0 70012 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_120_755
timestamp 1644511149
transform 1 0 70564 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_120_757
timestamp 1644511149
transform 1 0 70748 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_769
timestamp 1644511149
transform 1 0 71852 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_781
timestamp 1644511149
transform 1 0 72956 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_793
timestamp 1644511149
transform 1 0 74060 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_120_805
timestamp 1644511149
transform 1 0 75164 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_120_811
timestamp 1644511149
transform 1 0 75716 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_120_813
timestamp 1644511149
transform 1 0 75900 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_120_825
timestamp 1644511149
transform 1 0 77004 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_120_831
timestamp 1644511149
transform 1 0 77556 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_120_838
timestamp 1644511149
transform 1 0 78200 0 1 67456
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_121_3
timestamp 1644511149
transform 1 0 1380 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_15
timestamp 1644511149
transform 1 0 2484 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_27
timestamp 1644511149
transform 1 0 3588 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_39
timestamp 1644511149
transform 1 0 4692 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_121_51
timestamp 1644511149
transform 1 0 5796 0 -1 68544
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_121_55
timestamp 1644511149
transform 1 0 6164 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_121_57
timestamp 1644511149
transform 1 0 6348 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_69
timestamp 1644511149
transform 1 0 7452 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_81
timestamp 1644511149
transform 1 0 8556 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_93
timestamp 1644511149
transform 1 0 9660 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_121_105
timestamp 1644511149
transform 1 0 10764 0 -1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_121_111
timestamp 1644511149
transform 1 0 11316 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_121_113
timestamp 1644511149
transform 1 0 11500 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_125
timestamp 1644511149
transform 1 0 12604 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_137
timestamp 1644511149
transform 1 0 13708 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_149
timestamp 1644511149
transform 1 0 14812 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_121_161
timestamp 1644511149
transform 1 0 15916 0 -1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_121_167
timestamp 1644511149
transform 1 0 16468 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_121_169
timestamp 1644511149
transform 1 0 16652 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_181
timestamp 1644511149
transform 1 0 17756 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_193
timestamp 1644511149
transform 1 0 18860 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_205
timestamp 1644511149
transform 1 0 19964 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_121_217
timestamp 1644511149
transform 1 0 21068 0 -1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_121_223
timestamp 1644511149
transform 1 0 21620 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_121_225
timestamp 1644511149
transform 1 0 21804 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_237
timestamp 1644511149
transform 1 0 22908 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_249
timestamp 1644511149
transform 1 0 24012 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_261
timestamp 1644511149
transform 1 0 25116 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_121_273
timestamp 1644511149
transform 1 0 26220 0 -1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_121_279
timestamp 1644511149
transform 1 0 26772 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_121_281
timestamp 1644511149
transform 1 0 26956 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_293
timestamp 1644511149
transform 1 0 28060 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_305
timestamp 1644511149
transform 1 0 29164 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_317
timestamp 1644511149
transform 1 0 30268 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_121_329
timestamp 1644511149
transform 1 0 31372 0 -1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_121_335
timestamp 1644511149
transform 1 0 31924 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_121_337
timestamp 1644511149
transform 1 0 32108 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_349
timestamp 1644511149
transform 1 0 33212 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_361
timestamp 1644511149
transform 1 0 34316 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_373
timestamp 1644511149
transform 1 0 35420 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_121_385
timestamp 1644511149
transform 1 0 36524 0 -1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_121_391
timestamp 1644511149
transform 1 0 37076 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_121_393
timestamp 1644511149
transform 1 0 37260 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_405
timestamp 1644511149
transform 1 0 38364 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_417
timestamp 1644511149
transform 1 0 39468 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_429
timestamp 1644511149
transform 1 0 40572 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_121_441
timestamp 1644511149
transform 1 0 41676 0 -1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_121_447
timestamp 1644511149
transform 1 0 42228 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_121_449
timestamp 1644511149
transform 1 0 42412 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_461
timestamp 1644511149
transform 1 0 43516 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_473
timestamp 1644511149
transform 1 0 44620 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_485
timestamp 1644511149
transform 1 0 45724 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_121_497
timestamp 1644511149
transform 1 0 46828 0 -1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_121_503
timestamp 1644511149
transform 1 0 47380 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_121_505
timestamp 1644511149
transform 1 0 47564 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_517
timestamp 1644511149
transform 1 0 48668 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_529
timestamp 1644511149
transform 1 0 49772 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_541
timestamp 1644511149
transform 1 0 50876 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_121_553
timestamp 1644511149
transform 1 0 51980 0 -1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_121_559
timestamp 1644511149
transform 1 0 52532 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_121_561
timestamp 1644511149
transform 1 0 52716 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_573
timestamp 1644511149
transform 1 0 53820 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_585
timestamp 1644511149
transform 1 0 54924 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_597
timestamp 1644511149
transform 1 0 56028 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_121_609
timestamp 1644511149
transform 1 0 57132 0 -1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_121_615
timestamp 1644511149
transform 1 0 57684 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_121_617
timestamp 1644511149
transform 1 0 57868 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_629
timestamp 1644511149
transform 1 0 58972 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_641
timestamp 1644511149
transform 1 0 60076 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_653
timestamp 1644511149
transform 1 0 61180 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_121_665
timestamp 1644511149
transform 1 0 62284 0 -1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_121_671
timestamp 1644511149
transform 1 0 62836 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_121_673
timestamp 1644511149
transform 1 0 63020 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_685
timestamp 1644511149
transform 1 0 64124 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_697
timestamp 1644511149
transform 1 0 65228 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_709
timestamp 1644511149
transform 1 0 66332 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_121_721
timestamp 1644511149
transform 1 0 67436 0 -1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_121_727
timestamp 1644511149
transform 1 0 67988 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_121_729
timestamp 1644511149
transform 1 0 68172 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_741
timestamp 1644511149
transform 1 0 69276 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_753
timestamp 1644511149
transform 1 0 70380 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_765
timestamp 1644511149
transform 1 0 71484 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_121_777
timestamp 1644511149
transform 1 0 72588 0 -1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_121_783
timestamp 1644511149
transform 1 0 73140 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_121_785
timestamp 1644511149
transform 1 0 73324 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_797
timestamp 1644511149
transform 1 0 74428 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_809
timestamp 1644511149
transform 1 0 75532 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_821
timestamp 1644511149
transform 1 0 76636 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_121_833
timestamp 1644511149
transform 1 0 77740 0 -1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_121_839
timestamp 1644511149
transform 1 0 78292 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_121_841
timestamp 1644511149
transform 1 0 78476 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_122_3
timestamp 1644511149
transform 1 0 1380 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_15
timestamp 1644511149
transform 1 0 2484 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_122_27
timestamp 1644511149
transform 1 0 3588 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_122_29
timestamp 1644511149
transform 1 0 3772 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_41
timestamp 1644511149
transform 1 0 4876 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_53
timestamp 1644511149
transform 1 0 5980 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_65
timestamp 1644511149
transform 1 0 7084 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_122_77
timestamp 1644511149
transform 1 0 8188 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_122_83
timestamp 1644511149
transform 1 0 8740 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_122_85
timestamp 1644511149
transform 1 0 8924 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_97
timestamp 1644511149
transform 1 0 10028 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_109
timestamp 1644511149
transform 1 0 11132 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_121
timestamp 1644511149
transform 1 0 12236 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_122_133
timestamp 1644511149
transform 1 0 13340 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_122_139
timestamp 1644511149
transform 1 0 13892 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_122_141
timestamp 1644511149
transform 1 0 14076 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_153
timestamp 1644511149
transform 1 0 15180 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_165
timestamp 1644511149
transform 1 0 16284 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_177
timestamp 1644511149
transform 1 0 17388 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_122_189
timestamp 1644511149
transform 1 0 18492 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_122_195
timestamp 1644511149
transform 1 0 19044 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_122_197
timestamp 1644511149
transform 1 0 19228 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_209
timestamp 1644511149
transform 1 0 20332 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_221
timestamp 1644511149
transform 1 0 21436 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_233
timestamp 1644511149
transform 1 0 22540 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_122_245
timestamp 1644511149
transform 1 0 23644 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_122_251
timestamp 1644511149
transform 1 0 24196 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_122_253
timestamp 1644511149
transform 1 0 24380 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_265
timestamp 1644511149
transform 1 0 25484 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_277
timestamp 1644511149
transform 1 0 26588 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_289
timestamp 1644511149
transform 1 0 27692 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_122_301
timestamp 1644511149
transform 1 0 28796 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_122_307
timestamp 1644511149
transform 1 0 29348 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_122_309
timestamp 1644511149
transform 1 0 29532 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_321
timestamp 1644511149
transform 1 0 30636 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_333
timestamp 1644511149
transform 1 0 31740 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_345
timestamp 1644511149
transform 1 0 32844 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_122_357
timestamp 1644511149
transform 1 0 33948 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_122_363
timestamp 1644511149
transform 1 0 34500 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_122_365
timestamp 1644511149
transform 1 0 34684 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_377
timestamp 1644511149
transform 1 0 35788 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_389
timestamp 1644511149
transform 1 0 36892 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_401
timestamp 1644511149
transform 1 0 37996 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_122_413
timestamp 1644511149
transform 1 0 39100 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_122_419
timestamp 1644511149
transform 1 0 39652 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_122_421
timestamp 1644511149
transform 1 0 39836 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_433
timestamp 1644511149
transform 1 0 40940 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_445
timestamp 1644511149
transform 1 0 42044 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_457
timestamp 1644511149
transform 1 0 43148 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_122_469
timestamp 1644511149
transform 1 0 44252 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_122_475
timestamp 1644511149
transform 1 0 44804 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_122_477
timestamp 1644511149
transform 1 0 44988 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_489
timestamp 1644511149
transform 1 0 46092 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_501
timestamp 1644511149
transform 1 0 47196 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_513
timestamp 1644511149
transform 1 0 48300 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_122_525
timestamp 1644511149
transform 1 0 49404 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_122_531
timestamp 1644511149
transform 1 0 49956 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_122_533
timestamp 1644511149
transform 1 0 50140 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_545
timestamp 1644511149
transform 1 0 51244 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_557
timestamp 1644511149
transform 1 0 52348 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_569
timestamp 1644511149
transform 1 0 53452 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_122_581
timestamp 1644511149
transform 1 0 54556 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_122_587
timestamp 1644511149
transform 1 0 55108 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_122_589
timestamp 1644511149
transform 1 0 55292 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_601
timestamp 1644511149
transform 1 0 56396 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_613
timestamp 1644511149
transform 1 0 57500 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_625
timestamp 1644511149
transform 1 0 58604 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_122_637
timestamp 1644511149
transform 1 0 59708 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_122_643
timestamp 1644511149
transform 1 0 60260 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_122_645
timestamp 1644511149
transform 1 0 60444 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_657
timestamp 1644511149
transform 1 0 61548 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_669
timestamp 1644511149
transform 1 0 62652 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_681
timestamp 1644511149
transform 1 0 63756 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_122_693
timestamp 1644511149
transform 1 0 64860 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_122_699
timestamp 1644511149
transform 1 0 65412 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_122_701
timestamp 1644511149
transform 1 0 65596 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_713
timestamp 1644511149
transform 1 0 66700 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_725
timestamp 1644511149
transform 1 0 67804 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_737
timestamp 1644511149
transform 1 0 68908 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_122_749
timestamp 1644511149
transform 1 0 70012 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_122_755
timestamp 1644511149
transform 1 0 70564 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_122_757
timestamp 1644511149
transform 1 0 70748 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_769
timestamp 1644511149
transform 1 0 71852 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_781
timestamp 1644511149
transform 1 0 72956 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_793
timestamp 1644511149
transform 1 0 74060 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_122_805
timestamp 1644511149
transform 1 0 75164 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_122_811
timestamp 1644511149
transform 1 0 75716 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_122_813
timestamp 1644511149
transform 1 0 75900 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_825
timestamp 1644511149
transform 1 0 77004 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_122_837
timestamp 1644511149
transform 1 0 78108 0 1 68544
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_122_841
timestamp 1644511149
transform 1 0 78476 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_123_3
timestamp 1644511149
transform 1 0 1380 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_123_15
timestamp 1644511149
transform 1 0 2484 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_123_27
timestamp 1644511149
transform 1 0 3588 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_123_39
timestamp 1644511149
transform 1 0 4692 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_123_51
timestamp 1644511149
transform 1 0 5796 0 -1 69632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_123_55
timestamp 1644511149
transform 1 0 6164 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_123_57
timestamp 1644511149
transform 1 0 6348 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_123_69
timestamp 1644511149
transform 1 0 7452 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_123_81
timestamp 1644511149
transform 1 0 8556 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_123_93
timestamp 1644511149
transform 1 0 9660 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_123_105
timestamp 1644511149
transform 1 0 10764 0 -1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_123_111
timestamp 1644511149
transform 1 0 11316 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_123_113
timestamp 1644511149
transform 1 0 11500 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_123_125
timestamp 1644511149
transform 1 0 12604 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_123_137
timestamp 1644511149
transform 1 0 13708 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_123_149
timestamp 1644511149
transform 1 0 14812 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_123_161
timestamp 1644511149
transform 1 0 15916 0 -1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_123_167
timestamp 1644511149
transform 1 0 16468 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_123_169
timestamp 1644511149
transform 1 0 16652 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_123_181
timestamp 1644511149
transform 1 0 17756 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_123_193
timestamp 1644511149
transform 1 0 18860 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_123_205
timestamp 1644511149
transform 1 0 19964 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_123_217
timestamp 1644511149
transform 1 0 21068 0 -1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_123_223
timestamp 1644511149
transform 1 0 21620 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_123_225
timestamp 1644511149
transform 1 0 21804 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_123_237
timestamp 1644511149
transform 1 0 22908 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_123_249
timestamp 1644511149
transform 1 0 24012 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_123_261
timestamp 1644511149
transform 1 0 25116 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_123_273
timestamp 1644511149
transform 1 0 26220 0 -1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_123_279
timestamp 1644511149
transform 1 0 26772 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_123_281
timestamp 1644511149
transform 1 0 26956 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_123_293
timestamp 1644511149
transform 1 0 28060 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_123_305
timestamp 1644511149
transform 1 0 29164 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_123_317
timestamp 1644511149
transform 1 0 30268 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_123_329
timestamp 1644511149
transform 1 0 31372 0 -1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_123_335
timestamp 1644511149
transform 1 0 31924 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_123_337
timestamp 1644511149
transform 1 0 32108 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_123_349
timestamp 1644511149
transform 1 0 33212 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_123_361
timestamp 1644511149
transform 1 0 34316 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_123_373
timestamp 1644511149
transform 1 0 35420 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_123_385
timestamp 1644511149
transform 1 0 36524 0 -1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_123_391
timestamp 1644511149
transform 1 0 37076 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_123_393
timestamp 1644511149
transform 1 0 37260 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_123_405
timestamp 1644511149
transform 1 0 38364 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_123_417
timestamp 1644511149
transform 1 0 39468 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_123_429
timestamp 1644511149
transform 1 0 40572 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_123_441
timestamp 1644511149
transform 1 0 41676 0 -1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_123_447
timestamp 1644511149
transform 1 0 42228 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_123_449
timestamp 1644511149
transform 1 0 42412 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_123_461
timestamp 1644511149
transform 1 0 43516 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_123_473
timestamp 1644511149
transform 1 0 44620 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_123_485
timestamp 1644511149
transform 1 0 45724 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_123_497
timestamp 1644511149
transform 1 0 46828 0 -1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_123_503
timestamp 1644511149
transform 1 0 47380 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_123_505
timestamp 1644511149
transform 1 0 47564 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_123_517
timestamp 1644511149
transform 1 0 48668 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_123_529
timestamp 1644511149
transform 1 0 49772 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_123_541
timestamp 1644511149
transform 1 0 50876 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_123_553
timestamp 1644511149
transform 1 0 51980 0 -1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_123_559
timestamp 1644511149
transform 1 0 52532 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_123_561
timestamp 1644511149
transform 1 0 52716 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_123_573
timestamp 1644511149
transform 1 0 53820 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_123_585
timestamp 1644511149
transform 1 0 54924 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_123_597
timestamp 1644511149
transform 1 0 56028 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_123_609
timestamp 1644511149
transform 1 0 57132 0 -1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_123_615
timestamp 1644511149
transform 1 0 57684 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_123_617
timestamp 1644511149
transform 1 0 57868 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_123_629
timestamp 1644511149
transform 1 0 58972 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_123_641
timestamp 1644511149
transform 1 0 60076 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_123_653
timestamp 1644511149
transform 1 0 61180 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_123_665
timestamp 1644511149
transform 1 0 62284 0 -1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_123_671
timestamp 1644511149
transform 1 0 62836 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_123_673
timestamp 1644511149
transform 1 0 63020 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_123_685
timestamp 1644511149
transform 1 0 64124 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_123_697
timestamp 1644511149
transform 1 0 65228 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_123_709
timestamp 1644511149
transform 1 0 66332 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_123_721
timestamp 1644511149
transform 1 0 67436 0 -1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_123_727
timestamp 1644511149
transform 1 0 67988 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_123_729
timestamp 1644511149
transform 1 0 68172 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_123_741
timestamp 1644511149
transform 1 0 69276 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_123_753
timestamp 1644511149
transform 1 0 70380 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_123_765
timestamp 1644511149
transform 1 0 71484 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_123_777
timestamp 1644511149
transform 1 0 72588 0 -1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_123_783
timestamp 1644511149
transform 1 0 73140 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_123_785
timestamp 1644511149
transform 1 0 73324 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_123_797
timestamp 1644511149
transform 1 0 74428 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_123_809
timestamp 1644511149
transform 1 0 75532 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_123_821
timestamp 1644511149
transform 1 0 76636 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_123_833
timestamp 1644511149
transform 1 0 77740 0 -1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_123_839
timestamp 1644511149
transform 1 0 78292 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_123_841
timestamp 1644511149
transform 1 0 78476 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_124_3
timestamp 1644511149
transform 1 0 1380 0 1 69632
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_124_10
timestamp 1644511149
transform 1 0 2024 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_124_22
timestamp 1644511149
transform 1 0 3128 0 1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_124_29
timestamp 1644511149
transform 1 0 3772 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_124_41
timestamp 1644511149
transform 1 0 4876 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_124_53
timestamp 1644511149
transform 1 0 5980 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_124_65
timestamp 1644511149
transform 1 0 7084 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_124_77
timestamp 1644511149
transform 1 0 8188 0 1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_124_83
timestamp 1644511149
transform 1 0 8740 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_124_85
timestamp 1644511149
transform 1 0 8924 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_124_97
timestamp 1644511149
transform 1 0 10028 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_124_109
timestamp 1644511149
transform 1 0 11132 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_124_121
timestamp 1644511149
transform 1 0 12236 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_124_133
timestamp 1644511149
transform 1 0 13340 0 1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_124_139
timestamp 1644511149
transform 1 0 13892 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_124_141
timestamp 1644511149
transform 1 0 14076 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_124_153
timestamp 1644511149
transform 1 0 15180 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_124_165
timestamp 1644511149
transform 1 0 16284 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_124_177
timestamp 1644511149
transform 1 0 17388 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_124_189
timestamp 1644511149
transform 1 0 18492 0 1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_124_195
timestamp 1644511149
transform 1 0 19044 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_124_197
timestamp 1644511149
transform 1 0 19228 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_124_209
timestamp 1644511149
transform 1 0 20332 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_124_221
timestamp 1644511149
transform 1 0 21436 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_124_233
timestamp 1644511149
transform 1 0 22540 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_124_245
timestamp 1644511149
transform 1 0 23644 0 1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_124_251
timestamp 1644511149
transform 1 0 24196 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_124_253
timestamp 1644511149
transform 1 0 24380 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_124_265
timestamp 1644511149
transform 1 0 25484 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_124_277
timestamp 1644511149
transform 1 0 26588 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_124_289
timestamp 1644511149
transform 1 0 27692 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_124_301
timestamp 1644511149
transform 1 0 28796 0 1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_124_307
timestamp 1644511149
transform 1 0 29348 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_124_309
timestamp 1644511149
transform 1 0 29532 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_124_321
timestamp 1644511149
transform 1 0 30636 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_124_333
timestamp 1644511149
transform 1 0 31740 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_124_345
timestamp 1644511149
transform 1 0 32844 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_124_357
timestamp 1644511149
transform 1 0 33948 0 1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_124_363
timestamp 1644511149
transform 1 0 34500 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_124_365
timestamp 1644511149
transform 1 0 34684 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_124_377
timestamp 1644511149
transform 1 0 35788 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_124_389
timestamp 1644511149
transform 1 0 36892 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_124_401
timestamp 1644511149
transform 1 0 37996 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_124_413
timestamp 1644511149
transform 1 0 39100 0 1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_124_419
timestamp 1644511149
transform 1 0 39652 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_124_421
timestamp 1644511149
transform 1 0 39836 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_124_433
timestamp 1644511149
transform 1 0 40940 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_124_445
timestamp 1644511149
transform 1 0 42044 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_124_457
timestamp 1644511149
transform 1 0 43148 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_124_469
timestamp 1644511149
transform 1 0 44252 0 1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_124_475
timestamp 1644511149
transform 1 0 44804 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_124_477
timestamp 1644511149
transform 1 0 44988 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_124_489
timestamp 1644511149
transform 1 0 46092 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_124_501
timestamp 1644511149
transform 1 0 47196 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_124_513
timestamp 1644511149
transform 1 0 48300 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_124_525
timestamp 1644511149
transform 1 0 49404 0 1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_124_531
timestamp 1644511149
transform 1 0 49956 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_124_533
timestamp 1644511149
transform 1 0 50140 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_124_545
timestamp 1644511149
transform 1 0 51244 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_124_557
timestamp 1644511149
transform 1 0 52348 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_124_569
timestamp 1644511149
transform 1 0 53452 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_124_581
timestamp 1644511149
transform 1 0 54556 0 1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_124_587
timestamp 1644511149
transform 1 0 55108 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_124_589
timestamp 1644511149
transform 1 0 55292 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_124_601
timestamp 1644511149
transform 1 0 56396 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_124_613
timestamp 1644511149
transform 1 0 57500 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_124_625
timestamp 1644511149
transform 1 0 58604 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_124_637
timestamp 1644511149
transform 1 0 59708 0 1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_124_643
timestamp 1644511149
transform 1 0 60260 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_124_645
timestamp 1644511149
transform 1 0 60444 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_124_657
timestamp 1644511149
transform 1 0 61548 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_124_669
timestamp 1644511149
transform 1 0 62652 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_124_681
timestamp 1644511149
transform 1 0 63756 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_124_693
timestamp 1644511149
transform 1 0 64860 0 1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_124_699
timestamp 1644511149
transform 1 0 65412 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_124_701
timestamp 1644511149
transform 1 0 65596 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_124_713
timestamp 1644511149
transform 1 0 66700 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_124_725
timestamp 1644511149
transform 1 0 67804 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_124_737
timestamp 1644511149
transform 1 0 68908 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_124_749
timestamp 1644511149
transform 1 0 70012 0 1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_124_755
timestamp 1644511149
transform 1 0 70564 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_124_757
timestamp 1644511149
transform 1 0 70748 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_124_769
timestamp 1644511149
transform 1 0 71852 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_124_781
timestamp 1644511149
transform 1 0 72956 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_124_793
timestamp 1644511149
transform 1 0 74060 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_124_805
timestamp 1644511149
transform 1 0 75164 0 1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_124_811
timestamp 1644511149
transform 1 0 75716 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_124_813
timestamp 1644511149
transform 1 0 75900 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_124_825
timestamp 1644511149
transform 1 0 77004 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_124_837
timestamp 1644511149
transform 1 0 78108 0 1 69632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_124_841
timestamp 1644511149
transform 1 0 78476 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_125_7
timestamp 1644511149
transform 1 0 1748 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_125_19
timestamp 1644511149
transform 1 0 2852 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_125_31
timestamp 1644511149
transform 1 0 3956 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_125_43
timestamp 1644511149
transform 1 0 5060 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_125_55
timestamp 1644511149
transform 1 0 6164 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_125_57
timestamp 1644511149
transform 1 0 6348 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_125_69
timestamp 1644511149
transform 1 0 7452 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_125_81
timestamp 1644511149
transform 1 0 8556 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_125_93
timestamp 1644511149
transform 1 0 9660 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_125_105
timestamp 1644511149
transform 1 0 10764 0 -1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_125_111
timestamp 1644511149
transform 1 0 11316 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_125_113
timestamp 1644511149
transform 1 0 11500 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_125_125
timestamp 1644511149
transform 1 0 12604 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_125_137
timestamp 1644511149
transform 1 0 13708 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_125_149
timestamp 1644511149
transform 1 0 14812 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_125_161
timestamp 1644511149
transform 1 0 15916 0 -1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_125_167
timestamp 1644511149
transform 1 0 16468 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_125_169
timestamp 1644511149
transform 1 0 16652 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_125_181
timestamp 1644511149
transform 1 0 17756 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_125_193
timestamp 1644511149
transform 1 0 18860 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_125_205
timestamp 1644511149
transform 1 0 19964 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_125_217
timestamp 1644511149
transform 1 0 21068 0 -1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_125_223
timestamp 1644511149
transform 1 0 21620 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_125_225
timestamp 1644511149
transform 1 0 21804 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_125_237
timestamp 1644511149
transform 1 0 22908 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_125_249
timestamp 1644511149
transform 1 0 24012 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_125_261
timestamp 1644511149
transform 1 0 25116 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_125_273
timestamp 1644511149
transform 1 0 26220 0 -1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_125_279
timestamp 1644511149
transform 1 0 26772 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_125_281
timestamp 1644511149
transform 1 0 26956 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_125_293
timestamp 1644511149
transform 1 0 28060 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_125_305
timestamp 1644511149
transform 1 0 29164 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_125_317
timestamp 1644511149
transform 1 0 30268 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_125_329
timestamp 1644511149
transform 1 0 31372 0 -1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_125_335
timestamp 1644511149
transform 1 0 31924 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_125_337
timestamp 1644511149
transform 1 0 32108 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_125_349
timestamp 1644511149
transform 1 0 33212 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_125_361
timestamp 1644511149
transform 1 0 34316 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_125_373
timestamp 1644511149
transform 1 0 35420 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_125_385
timestamp 1644511149
transform 1 0 36524 0 -1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_125_391
timestamp 1644511149
transform 1 0 37076 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_125_393
timestamp 1644511149
transform 1 0 37260 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_125_405
timestamp 1644511149
transform 1 0 38364 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_125_417
timestamp 1644511149
transform 1 0 39468 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_125_429
timestamp 1644511149
transform 1 0 40572 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_125_441
timestamp 1644511149
transform 1 0 41676 0 -1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_125_447
timestamp 1644511149
transform 1 0 42228 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_125_449
timestamp 1644511149
transform 1 0 42412 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_125_461
timestamp 1644511149
transform 1 0 43516 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_125_473
timestamp 1644511149
transform 1 0 44620 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_125_485
timestamp 1644511149
transform 1 0 45724 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_125_497
timestamp 1644511149
transform 1 0 46828 0 -1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_125_503
timestamp 1644511149
transform 1 0 47380 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_125_505
timestamp 1644511149
transform 1 0 47564 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_125_517
timestamp 1644511149
transform 1 0 48668 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_125_529
timestamp 1644511149
transform 1 0 49772 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_125_541
timestamp 1644511149
transform 1 0 50876 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_125_553
timestamp 1644511149
transform 1 0 51980 0 -1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_125_559
timestamp 1644511149
transform 1 0 52532 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_125_561
timestamp 1644511149
transform 1 0 52716 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_125_573
timestamp 1644511149
transform 1 0 53820 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_125_585
timestamp 1644511149
transform 1 0 54924 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_125_597
timestamp 1644511149
transform 1 0 56028 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_125_609
timestamp 1644511149
transform 1 0 57132 0 -1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_125_615
timestamp 1644511149
transform 1 0 57684 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_125_617
timestamp 1644511149
transform 1 0 57868 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_125_629
timestamp 1644511149
transform 1 0 58972 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_125_641
timestamp 1644511149
transform 1 0 60076 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_125_653
timestamp 1644511149
transform 1 0 61180 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_125_665
timestamp 1644511149
transform 1 0 62284 0 -1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_125_671
timestamp 1644511149
transform 1 0 62836 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_125_673
timestamp 1644511149
transform 1 0 63020 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_125_685
timestamp 1644511149
transform 1 0 64124 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_125_697
timestamp 1644511149
transform 1 0 65228 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_125_709
timestamp 1644511149
transform 1 0 66332 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_125_721
timestamp 1644511149
transform 1 0 67436 0 -1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_125_727
timestamp 1644511149
transform 1 0 67988 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_125_729
timestamp 1644511149
transform 1 0 68172 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_125_741
timestamp 1644511149
transform 1 0 69276 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_125_753
timestamp 1644511149
transform 1 0 70380 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_125_765
timestamp 1644511149
transform 1 0 71484 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_125_777
timestamp 1644511149
transform 1 0 72588 0 -1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_125_783
timestamp 1644511149
transform 1 0 73140 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_125_785
timestamp 1644511149
transform 1 0 73324 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_125_797
timestamp 1644511149
transform 1 0 74428 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_125_809
timestamp 1644511149
transform 1 0 75532 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_125_821
timestamp 1644511149
transform 1 0 76636 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_125_833
timestamp 1644511149
transform 1 0 77740 0 -1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_125_839
timestamp 1644511149
transform 1 0 78292 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_125_841
timestamp 1644511149
transform 1 0 78476 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_126_3
timestamp 1644511149
transform 1 0 1380 0 1 70720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_126_11
timestamp 1644511149
transform 1 0 2116 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_126_23
timestamp 1644511149
transform 1 0 3220 0 1 70720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_126_27
timestamp 1644511149
transform 1 0 3588 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_126_29
timestamp 1644511149
transform 1 0 3772 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_126_41
timestamp 1644511149
transform 1 0 4876 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_126_53
timestamp 1644511149
transform 1 0 5980 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_126_65
timestamp 1644511149
transform 1 0 7084 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_126_77
timestamp 1644511149
transform 1 0 8188 0 1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_126_83
timestamp 1644511149
transform 1 0 8740 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_126_85
timestamp 1644511149
transform 1 0 8924 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_126_97
timestamp 1644511149
transform 1 0 10028 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_126_109
timestamp 1644511149
transform 1 0 11132 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_126_121
timestamp 1644511149
transform 1 0 12236 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_126_133
timestamp 1644511149
transform 1 0 13340 0 1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_126_139
timestamp 1644511149
transform 1 0 13892 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_126_141
timestamp 1644511149
transform 1 0 14076 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_126_153
timestamp 1644511149
transform 1 0 15180 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_126_165
timestamp 1644511149
transform 1 0 16284 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_126_177
timestamp 1644511149
transform 1 0 17388 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_126_189
timestamp 1644511149
transform 1 0 18492 0 1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_126_195
timestamp 1644511149
transform 1 0 19044 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_126_197
timestamp 1644511149
transform 1 0 19228 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_126_209
timestamp 1644511149
transform 1 0 20332 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_126_221
timestamp 1644511149
transform 1 0 21436 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_126_233
timestamp 1644511149
transform 1 0 22540 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_126_245
timestamp 1644511149
transform 1 0 23644 0 1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_126_251
timestamp 1644511149
transform 1 0 24196 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_126_253
timestamp 1644511149
transform 1 0 24380 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_126_265
timestamp 1644511149
transform 1 0 25484 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_126_277
timestamp 1644511149
transform 1 0 26588 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_126_289
timestamp 1644511149
transform 1 0 27692 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_126_301
timestamp 1644511149
transform 1 0 28796 0 1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_126_307
timestamp 1644511149
transform 1 0 29348 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_126_309
timestamp 1644511149
transform 1 0 29532 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_126_321
timestamp 1644511149
transform 1 0 30636 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_126_333
timestamp 1644511149
transform 1 0 31740 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_126_345
timestamp 1644511149
transform 1 0 32844 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_126_357
timestamp 1644511149
transform 1 0 33948 0 1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_126_363
timestamp 1644511149
transform 1 0 34500 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_126_365
timestamp 1644511149
transform 1 0 34684 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_126_377
timestamp 1644511149
transform 1 0 35788 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_126_389
timestamp 1644511149
transform 1 0 36892 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_126_401
timestamp 1644511149
transform 1 0 37996 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_126_413
timestamp 1644511149
transform 1 0 39100 0 1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_126_419
timestamp 1644511149
transform 1 0 39652 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_126_421
timestamp 1644511149
transform 1 0 39836 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_126_433
timestamp 1644511149
transform 1 0 40940 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_126_445
timestamp 1644511149
transform 1 0 42044 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_126_457
timestamp 1644511149
transform 1 0 43148 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_126_469
timestamp 1644511149
transform 1 0 44252 0 1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_126_475
timestamp 1644511149
transform 1 0 44804 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_126_477
timestamp 1644511149
transform 1 0 44988 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_126_489
timestamp 1644511149
transform 1 0 46092 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_126_501
timestamp 1644511149
transform 1 0 47196 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_126_513
timestamp 1644511149
transform 1 0 48300 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_126_525
timestamp 1644511149
transform 1 0 49404 0 1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_126_531
timestamp 1644511149
transform 1 0 49956 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_126_533
timestamp 1644511149
transform 1 0 50140 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_126_545
timestamp 1644511149
transform 1 0 51244 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_126_557
timestamp 1644511149
transform 1 0 52348 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_126_569
timestamp 1644511149
transform 1 0 53452 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_126_581
timestamp 1644511149
transform 1 0 54556 0 1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_126_587
timestamp 1644511149
transform 1 0 55108 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_126_589
timestamp 1644511149
transform 1 0 55292 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_126_601
timestamp 1644511149
transform 1 0 56396 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_126_613
timestamp 1644511149
transform 1 0 57500 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_126_625
timestamp 1644511149
transform 1 0 58604 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_126_637
timestamp 1644511149
transform 1 0 59708 0 1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_126_643
timestamp 1644511149
transform 1 0 60260 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_126_645
timestamp 1644511149
transform 1 0 60444 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_126_657
timestamp 1644511149
transform 1 0 61548 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_126_669
timestamp 1644511149
transform 1 0 62652 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_126_681
timestamp 1644511149
transform 1 0 63756 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_126_693
timestamp 1644511149
transform 1 0 64860 0 1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_126_699
timestamp 1644511149
transform 1 0 65412 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_126_701
timestamp 1644511149
transform 1 0 65596 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_126_713
timestamp 1644511149
transform 1 0 66700 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_126_725
timestamp 1644511149
transform 1 0 67804 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_126_737
timestamp 1644511149
transform 1 0 68908 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_126_749
timestamp 1644511149
transform 1 0 70012 0 1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_126_755
timestamp 1644511149
transform 1 0 70564 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_126_757
timestamp 1644511149
transform 1 0 70748 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_126_769
timestamp 1644511149
transform 1 0 71852 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_126_781
timestamp 1644511149
transform 1 0 72956 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_126_793
timestamp 1644511149
transform 1 0 74060 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_126_805
timestamp 1644511149
transform 1 0 75164 0 1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_126_811
timestamp 1644511149
transform 1 0 75716 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_126_813
timestamp 1644511149
transform 1 0 75900 0 1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_126_819
timestamp 1644511149
transform 1 0 76452 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_126_823
timestamp 1644511149
transform 1 0 76820 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_126_835
timestamp 1644511149
transform 1 0 77924 0 1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_126_841
timestamp 1644511149
transform 1 0 78476 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_127_3
timestamp 1644511149
transform 1 0 1380 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_127_15
timestamp 1644511149
transform 1 0 2484 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_127_27
timestamp 1644511149
transform 1 0 3588 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_127_39
timestamp 1644511149
transform 1 0 4692 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_127_51
timestamp 1644511149
transform 1 0 5796 0 -1 71808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_127_55
timestamp 1644511149
transform 1 0 6164 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_127_57
timestamp 1644511149
transform 1 0 6348 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_127_69
timestamp 1644511149
transform 1 0 7452 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_127_81
timestamp 1644511149
transform 1 0 8556 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_127_93
timestamp 1644511149
transform 1 0 9660 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_127_105
timestamp 1644511149
transform 1 0 10764 0 -1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_127_111
timestamp 1644511149
transform 1 0 11316 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_127_113
timestamp 1644511149
transform 1 0 11500 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_127_125
timestamp 1644511149
transform 1 0 12604 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_127_137
timestamp 1644511149
transform 1 0 13708 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_127_149
timestamp 1644511149
transform 1 0 14812 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_127_161
timestamp 1644511149
transform 1 0 15916 0 -1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_127_167
timestamp 1644511149
transform 1 0 16468 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_127_169
timestamp 1644511149
transform 1 0 16652 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_127_181
timestamp 1644511149
transform 1 0 17756 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_127_193
timestamp 1644511149
transform 1 0 18860 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_127_205
timestamp 1644511149
transform 1 0 19964 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_127_217
timestamp 1644511149
transform 1 0 21068 0 -1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_127_223
timestamp 1644511149
transform 1 0 21620 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_127_225
timestamp 1644511149
transform 1 0 21804 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_127_237
timestamp 1644511149
transform 1 0 22908 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_127_249
timestamp 1644511149
transform 1 0 24012 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_127_261
timestamp 1644511149
transform 1 0 25116 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_127_273
timestamp 1644511149
transform 1 0 26220 0 -1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_127_279
timestamp 1644511149
transform 1 0 26772 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_127_281
timestamp 1644511149
transform 1 0 26956 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_127_293
timestamp 1644511149
transform 1 0 28060 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_127_305
timestamp 1644511149
transform 1 0 29164 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_127_317
timestamp 1644511149
transform 1 0 30268 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_127_329
timestamp 1644511149
transform 1 0 31372 0 -1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_127_335
timestamp 1644511149
transform 1 0 31924 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_127_337
timestamp 1644511149
transform 1 0 32108 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_127_349
timestamp 1644511149
transform 1 0 33212 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_127_361
timestamp 1644511149
transform 1 0 34316 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_127_373
timestamp 1644511149
transform 1 0 35420 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_127_385
timestamp 1644511149
transform 1 0 36524 0 -1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_127_391
timestamp 1644511149
transform 1 0 37076 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_127_393
timestamp 1644511149
transform 1 0 37260 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_127_405
timestamp 1644511149
transform 1 0 38364 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_127_417
timestamp 1644511149
transform 1 0 39468 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_127_429
timestamp 1644511149
transform 1 0 40572 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_127_441
timestamp 1644511149
transform 1 0 41676 0 -1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_127_447
timestamp 1644511149
transform 1 0 42228 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_127_449
timestamp 1644511149
transform 1 0 42412 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_127_461
timestamp 1644511149
transform 1 0 43516 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_127_473
timestamp 1644511149
transform 1 0 44620 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_127_485
timestamp 1644511149
transform 1 0 45724 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_127_497
timestamp 1644511149
transform 1 0 46828 0 -1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_127_503
timestamp 1644511149
transform 1 0 47380 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_127_505
timestamp 1644511149
transform 1 0 47564 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_127_517
timestamp 1644511149
transform 1 0 48668 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_127_529
timestamp 1644511149
transform 1 0 49772 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_127_541
timestamp 1644511149
transform 1 0 50876 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_127_553
timestamp 1644511149
transform 1 0 51980 0 -1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_127_559
timestamp 1644511149
transform 1 0 52532 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_127_561
timestamp 1644511149
transform 1 0 52716 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_127_573
timestamp 1644511149
transform 1 0 53820 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_127_585
timestamp 1644511149
transform 1 0 54924 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_127_597
timestamp 1644511149
transform 1 0 56028 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_127_609
timestamp 1644511149
transform 1 0 57132 0 -1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_127_615
timestamp 1644511149
transform 1 0 57684 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_127_617
timestamp 1644511149
transform 1 0 57868 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_127_629
timestamp 1644511149
transform 1 0 58972 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_127_641
timestamp 1644511149
transform 1 0 60076 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_127_653
timestamp 1644511149
transform 1 0 61180 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_127_665
timestamp 1644511149
transform 1 0 62284 0 -1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_127_671
timestamp 1644511149
transform 1 0 62836 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_127_673
timestamp 1644511149
transform 1 0 63020 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_127_685
timestamp 1644511149
transform 1 0 64124 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_127_697
timestamp 1644511149
transform 1 0 65228 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_127_709
timestamp 1644511149
transform 1 0 66332 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_127_721
timestamp 1644511149
transform 1 0 67436 0 -1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_127_727
timestamp 1644511149
transform 1 0 67988 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_127_729
timestamp 1644511149
transform 1 0 68172 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_127_741
timestamp 1644511149
transform 1 0 69276 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_127_753
timestamp 1644511149
transform 1 0 70380 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_127_765
timestamp 1644511149
transform 1 0 71484 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_127_777
timestamp 1644511149
transform 1 0 72588 0 -1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_127_783
timestamp 1644511149
transform 1 0 73140 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_127_785
timestamp 1644511149
transform 1 0 73324 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_127_797
timestamp 1644511149
transform 1 0 74428 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_127_809
timestamp 1644511149
transform 1 0 75532 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_127_821
timestamp 1644511149
transform 1 0 76636 0 -1 71808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_127_829
timestamp 1644511149
transform 1 0 77372 0 -1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_127_836
timestamp 1644511149
transform 1 0 78016 0 -1 71808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_127_841
timestamp 1644511149
transform 1 0 78476 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_128_3
timestamp 1644511149
transform 1 0 1380 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_128_15
timestamp 1644511149
transform 1 0 2484 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_128_27
timestamp 1644511149
transform 1 0 3588 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_128_29
timestamp 1644511149
transform 1 0 3772 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_128_41
timestamp 1644511149
transform 1 0 4876 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_128_53
timestamp 1644511149
transform 1 0 5980 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_128_65
timestamp 1644511149
transform 1 0 7084 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_128_77
timestamp 1644511149
transform 1 0 8188 0 1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_128_83
timestamp 1644511149
transform 1 0 8740 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_128_85
timestamp 1644511149
transform 1 0 8924 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_128_97
timestamp 1644511149
transform 1 0 10028 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_128_109
timestamp 1644511149
transform 1 0 11132 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_128_121
timestamp 1644511149
transform 1 0 12236 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_128_133
timestamp 1644511149
transform 1 0 13340 0 1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_128_139
timestamp 1644511149
transform 1 0 13892 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_128_141
timestamp 1644511149
transform 1 0 14076 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_128_153
timestamp 1644511149
transform 1 0 15180 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_128_165
timestamp 1644511149
transform 1 0 16284 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_128_177
timestamp 1644511149
transform 1 0 17388 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_128_189
timestamp 1644511149
transform 1 0 18492 0 1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_128_195
timestamp 1644511149
transform 1 0 19044 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_128_197
timestamp 1644511149
transform 1 0 19228 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_128_209
timestamp 1644511149
transform 1 0 20332 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_128_221
timestamp 1644511149
transform 1 0 21436 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_128_233
timestamp 1644511149
transform 1 0 22540 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_128_245
timestamp 1644511149
transform 1 0 23644 0 1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_128_251
timestamp 1644511149
transform 1 0 24196 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_128_253
timestamp 1644511149
transform 1 0 24380 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_128_265
timestamp 1644511149
transform 1 0 25484 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_128_277
timestamp 1644511149
transform 1 0 26588 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_128_289
timestamp 1644511149
transform 1 0 27692 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_128_301
timestamp 1644511149
transform 1 0 28796 0 1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_128_307
timestamp 1644511149
transform 1 0 29348 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_128_309
timestamp 1644511149
transform 1 0 29532 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_128_321
timestamp 1644511149
transform 1 0 30636 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_128_333
timestamp 1644511149
transform 1 0 31740 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_128_345
timestamp 1644511149
transform 1 0 32844 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_128_357
timestamp 1644511149
transform 1 0 33948 0 1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_128_363
timestamp 1644511149
transform 1 0 34500 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_128_365
timestamp 1644511149
transform 1 0 34684 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_128_377
timestamp 1644511149
transform 1 0 35788 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_128_389
timestamp 1644511149
transform 1 0 36892 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_128_401
timestamp 1644511149
transform 1 0 37996 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_128_413
timestamp 1644511149
transform 1 0 39100 0 1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_128_419
timestamp 1644511149
transform 1 0 39652 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_128_421
timestamp 1644511149
transform 1 0 39836 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_128_433
timestamp 1644511149
transform 1 0 40940 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_128_445
timestamp 1644511149
transform 1 0 42044 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_128_457
timestamp 1644511149
transform 1 0 43148 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_128_469
timestamp 1644511149
transform 1 0 44252 0 1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_128_475
timestamp 1644511149
transform 1 0 44804 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_128_477
timestamp 1644511149
transform 1 0 44988 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_128_489
timestamp 1644511149
transform 1 0 46092 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_128_501
timestamp 1644511149
transform 1 0 47196 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_128_513
timestamp 1644511149
transform 1 0 48300 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_128_525
timestamp 1644511149
transform 1 0 49404 0 1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_128_531
timestamp 1644511149
transform 1 0 49956 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_128_533
timestamp 1644511149
transform 1 0 50140 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_128_545
timestamp 1644511149
transform 1 0 51244 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_128_557
timestamp 1644511149
transform 1 0 52348 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_128_569
timestamp 1644511149
transform 1 0 53452 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_128_581
timestamp 1644511149
transform 1 0 54556 0 1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_128_587
timestamp 1644511149
transform 1 0 55108 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_128_589
timestamp 1644511149
transform 1 0 55292 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_128_601
timestamp 1644511149
transform 1 0 56396 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_128_613
timestamp 1644511149
transform 1 0 57500 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_128_625
timestamp 1644511149
transform 1 0 58604 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_128_637
timestamp 1644511149
transform 1 0 59708 0 1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_128_643
timestamp 1644511149
transform 1 0 60260 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_128_645
timestamp 1644511149
transform 1 0 60444 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_128_657
timestamp 1644511149
transform 1 0 61548 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_128_669
timestamp 1644511149
transform 1 0 62652 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_128_681
timestamp 1644511149
transform 1 0 63756 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_128_693
timestamp 1644511149
transform 1 0 64860 0 1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_128_699
timestamp 1644511149
transform 1 0 65412 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_128_701
timestamp 1644511149
transform 1 0 65596 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_128_713
timestamp 1644511149
transform 1 0 66700 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_128_731
timestamp 1644511149
transform 1 0 68356 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_128_743
timestamp 1644511149
transform 1 0 69460 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_128_755
timestamp 1644511149
transform 1 0 70564 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_128_757
timestamp 1644511149
transform 1 0 70748 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_128_769
timestamp 1644511149
transform 1 0 71852 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_128_781
timestamp 1644511149
transform 1 0 72956 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_128_793
timestamp 1644511149
transform 1 0 74060 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_128_805
timestamp 1644511149
transform 1 0 75164 0 1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_128_811
timestamp 1644511149
transform 1 0 75716 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_128_813
timestamp 1644511149
transform 1 0 75900 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_128_825
timestamp 1644511149
transform 1 0 77004 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_128_837
timestamp 1644511149
transform 1 0 78108 0 1 71808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_128_841
timestamp 1644511149
transform 1 0 78476 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_129_3
timestamp 1644511149
transform 1 0 1380 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_129_15
timestamp 1644511149
transform 1 0 2484 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_129_27
timestamp 1644511149
transform 1 0 3588 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_129_39
timestamp 1644511149
transform 1 0 4692 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_129_51
timestamp 1644511149
transform 1 0 5796 0 -1 72896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_129_55
timestamp 1644511149
transform 1 0 6164 0 -1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_129_57
timestamp 1644511149
transform 1 0 6348 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_129_69
timestamp 1644511149
transform 1 0 7452 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_129_81
timestamp 1644511149
transform 1 0 8556 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_129_93
timestamp 1644511149
transform 1 0 9660 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_129_105
timestamp 1644511149
transform 1 0 10764 0 -1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_129_111
timestamp 1644511149
transform 1 0 11316 0 -1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_129_113
timestamp 1644511149
transform 1 0 11500 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_129_125
timestamp 1644511149
transform 1 0 12604 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_129_137
timestamp 1644511149
transform 1 0 13708 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_129_149
timestamp 1644511149
transform 1 0 14812 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_129_161
timestamp 1644511149
transform 1 0 15916 0 -1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_129_167
timestamp 1644511149
transform 1 0 16468 0 -1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_129_169
timestamp 1644511149
transform 1 0 16652 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_129_181
timestamp 1644511149
transform 1 0 17756 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_129_193
timestamp 1644511149
transform 1 0 18860 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_129_205
timestamp 1644511149
transform 1 0 19964 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_129_217
timestamp 1644511149
transform 1 0 21068 0 -1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_129_223
timestamp 1644511149
transform 1 0 21620 0 -1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_129_225
timestamp 1644511149
transform 1 0 21804 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_129_237
timestamp 1644511149
transform 1 0 22908 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_129_249
timestamp 1644511149
transform 1 0 24012 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_129_261
timestamp 1644511149
transform 1 0 25116 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_129_273
timestamp 1644511149
transform 1 0 26220 0 -1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_129_279
timestamp 1644511149
transform 1 0 26772 0 -1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_129_281
timestamp 1644511149
transform 1 0 26956 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_129_293
timestamp 1644511149
transform 1 0 28060 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_129_305
timestamp 1644511149
transform 1 0 29164 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_129_317
timestamp 1644511149
transform 1 0 30268 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_129_329
timestamp 1644511149
transform 1 0 31372 0 -1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_129_335
timestamp 1644511149
transform 1 0 31924 0 -1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_129_337
timestamp 1644511149
transform 1 0 32108 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_129_349
timestamp 1644511149
transform 1 0 33212 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_129_361
timestamp 1644511149
transform 1 0 34316 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_129_373
timestamp 1644511149
transform 1 0 35420 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_129_385
timestamp 1644511149
transform 1 0 36524 0 -1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_129_391
timestamp 1644511149
transform 1 0 37076 0 -1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_129_393
timestamp 1644511149
transform 1 0 37260 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_129_405
timestamp 1644511149
transform 1 0 38364 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_129_417
timestamp 1644511149
transform 1 0 39468 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_129_429
timestamp 1644511149
transform 1 0 40572 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_129_441
timestamp 1644511149
transform 1 0 41676 0 -1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_129_447
timestamp 1644511149
transform 1 0 42228 0 -1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_129_449
timestamp 1644511149
transform 1 0 42412 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_129_461
timestamp 1644511149
transform 1 0 43516 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_129_473
timestamp 1644511149
transform 1 0 44620 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_129_485
timestamp 1644511149
transform 1 0 45724 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_129_497
timestamp 1644511149
transform 1 0 46828 0 -1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_129_503
timestamp 1644511149
transform 1 0 47380 0 -1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_129_505
timestamp 1644511149
transform 1 0 47564 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_129_517
timestamp 1644511149
transform 1 0 48668 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_129_529
timestamp 1644511149
transform 1 0 49772 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_129_541
timestamp 1644511149
transform 1 0 50876 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_129_553
timestamp 1644511149
transform 1 0 51980 0 -1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_129_559
timestamp 1644511149
transform 1 0 52532 0 -1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_129_561
timestamp 1644511149
transform 1 0 52716 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_129_573
timestamp 1644511149
transform 1 0 53820 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_129_585
timestamp 1644511149
transform 1 0 54924 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_129_597
timestamp 1644511149
transform 1 0 56028 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_129_609
timestamp 1644511149
transform 1 0 57132 0 -1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_129_615
timestamp 1644511149
transform 1 0 57684 0 -1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_129_617
timestamp 1644511149
transform 1 0 57868 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_129_629
timestamp 1644511149
transform 1 0 58972 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_129_641
timestamp 1644511149
transform 1 0 60076 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_129_653
timestamp 1644511149
transform 1 0 61180 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_129_665
timestamp 1644511149
transform 1 0 62284 0 -1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_129_671
timestamp 1644511149
transform 1 0 62836 0 -1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_129_673
timestamp 1644511149
transform 1 0 63020 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_129_685
timestamp 1644511149
transform 1 0 64124 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_129_697
timestamp 1644511149
transform 1 0 65228 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_129_709
timestamp 1644511149
transform 1 0 66332 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_129_721
timestamp 1644511149
transform 1 0 67436 0 -1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_129_727
timestamp 1644511149
transform 1 0 67988 0 -1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_129_729
timestamp 1644511149
transform 1 0 68172 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_129_741
timestamp 1644511149
transform 1 0 69276 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_129_753
timestamp 1644511149
transform 1 0 70380 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_129_765
timestamp 1644511149
transform 1 0 71484 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_129_777
timestamp 1644511149
transform 1 0 72588 0 -1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_129_783
timestamp 1644511149
transform 1 0 73140 0 -1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_129_785
timestamp 1644511149
transform 1 0 73324 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_129_797
timestamp 1644511149
transform 1 0 74428 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_129_809
timestamp 1644511149
transform 1 0 75532 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_129_821
timestamp 1644511149
transform 1 0 76636 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_129_833
timestamp 1644511149
transform 1 0 77740 0 -1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_129_839
timestamp 1644511149
transform 1 0 78292 0 -1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_129_841
timestamp 1644511149
transform 1 0 78476 0 -1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_130_3
timestamp 1644511149
transform 1 0 1380 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_130_15
timestamp 1644511149
transform 1 0 2484 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_130_27
timestamp 1644511149
transform 1 0 3588 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_130_29
timestamp 1644511149
transform 1 0 3772 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_130_41
timestamp 1644511149
transform 1 0 4876 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_130_53
timestamp 1644511149
transform 1 0 5980 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_130_65
timestamp 1644511149
transform 1 0 7084 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_130_77
timestamp 1644511149
transform 1 0 8188 0 1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_130_83
timestamp 1644511149
transform 1 0 8740 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_130_85
timestamp 1644511149
transform 1 0 8924 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_130_97
timestamp 1644511149
transform 1 0 10028 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_130_109
timestamp 1644511149
transform 1 0 11132 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_130_121
timestamp 1644511149
transform 1 0 12236 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_130_133
timestamp 1644511149
transform 1 0 13340 0 1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_130_139
timestamp 1644511149
transform 1 0 13892 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_130_141
timestamp 1644511149
transform 1 0 14076 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_130_153
timestamp 1644511149
transform 1 0 15180 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_130_165
timestamp 1644511149
transform 1 0 16284 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_130_177
timestamp 1644511149
transform 1 0 17388 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_130_189
timestamp 1644511149
transform 1 0 18492 0 1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_130_195
timestamp 1644511149
transform 1 0 19044 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_130_197
timestamp 1644511149
transform 1 0 19228 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_130_209
timestamp 1644511149
transform 1 0 20332 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_130_221
timestamp 1644511149
transform 1 0 21436 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_130_233
timestamp 1644511149
transform 1 0 22540 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_130_245
timestamp 1644511149
transform 1 0 23644 0 1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_130_251
timestamp 1644511149
transform 1 0 24196 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_130_253
timestamp 1644511149
transform 1 0 24380 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_130_265
timestamp 1644511149
transform 1 0 25484 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_130_277
timestamp 1644511149
transform 1 0 26588 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_130_289
timestamp 1644511149
transform 1 0 27692 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_130_301
timestamp 1644511149
transform 1 0 28796 0 1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_130_307
timestamp 1644511149
transform 1 0 29348 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_130_309
timestamp 1644511149
transform 1 0 29532 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_130_321
timestamp 1644511149
transform 1 0 30636 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_130_333
timestamp 1644511149
transform 1 0 31740 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_130_345
timestamp 1644511149
transform 1 0 32844 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_130_357
timestamp 1644511149
transform 1 0 33948 0 1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_130_363
timestamp 1644511149
transform 1 0 34500 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_130_365
timestamp 1644511149
transform 1 0 34684 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_130_377
timestamp 1644511149
transform 1 0 35788 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_130_389
timestamp 1644511149
transform 1 0 36892 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_130_401
timestamp 1644511149
transform 1 0 37996 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_130_413
timestamp 1644511149
transform 1 0 39100 0 1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_130_419
timestamp 1644511149
transform 1 0 39652 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_130_421
timestamp 1644511149
transform 1 0 39836 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_130_433
timestamp 1644511149
transform 1 0 40940 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_130_445
timestamp 1644511149
transform 1 0 42044 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_130_457
timestamp 1644511149
transform 1 0 43148 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_130_469
timestamp 1644511149
transform 1 0 44252 0 1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_130_475
timestamp 1644511149
transform 1 0 44804 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_130_477
timestamp 1644511149
transform 1 0 44988 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_130_489
timestamp 1644511149
transform 1 0 46092 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_130_501
timestamp 1644511149
transform 1 0 47196 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_130_513
timestamp 1644511149
transform 1 0 48300 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_130_525
timestamp 1644511149
transform 1 0 49404 0 1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_130_531
timestamp 1644511149
transform 1 0 49956 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_130_533
timestamp 1644511149
transform 1 0 50140 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_130_545
timestamp 1644511149
transform 1 0 51244 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_130_557
timestamp 1644511149
transform 1 0 52348 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_130_569
timestamp 1644511149
transform 1 0 53452 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_130_581
timestamp 1644511149
transform 1 0 54556 0 1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_130_587
timestamp 1644511149
transform 1 0 55108 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_130_589
timestamp 1644511149
transform 1 0 55292 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_130_601
timestamp 1644511149
transform 1 0 56396 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_130_613
timestamp 1644511149
transform 1 0 57500 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_130_625
timestamp 1644511149
transform 1 0 58604 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_130_637
timestamp 1644511149
transform 1 0 59708 0 1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_130_643
timestamp 1644511149
transform 1 0 60260 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_130_645
timestamp 1644511149
transform 1 0 60444 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_130_657
timestamp 1644511149
transform 1 0 61548 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_130_669
timestamp 1644511149
transform 1 0 62652 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_130_681
timestamp 1644511149
transform 1 0 63756 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_130_693
timestamp 1644511149
transform 1 0 64860 0 1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_130_699
timestamp 1644511149
transform 1 0 65412 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_130_701
timestamp 1644511149
transform 1 0 65596 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_130_713
timestamp 1644511149
transform 1 0 66700 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_130_725
timestamp 1644511149
transform 1 0 67804 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_130_737
timestamp 1644511149
transform 1 0 68908 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_130_749
timestamp 1644511149
transform 1 0 70012 0 1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_130_755
timestamp 1644511149
transform 1 0 70564 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_130_757
timestamp 1644511149
transform 1 0 70748 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_130_769
timestamp 1644511149
transform 1 0 71852 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_130_781
timestamp 1644511149
transform 1 0 72956 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_130_793
timestamp 1644511149
transform 1 0 74060 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_130_805
timestamp 1644511149
transform 1 0 75164 0 1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_130_811
timestamp 1644511149
transform 1 0 75716 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_130_813
timestamp 1644511149
transform 1 0 75900 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_130_825
timestamp 1644511149
transform 1 0 77004 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_130_837
timestamp 1644511149
transform 1 0 78108 0 1 72896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_130_841
timestamp 1644511149
transform 1 0 78476 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_131_3
timestamp 1644511149
transform 1 0 1380 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_131_15
timestamp 1644511149
transform 1 0 2484 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_131_27
timestamp 1644511149
transform 1 0 3588 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_131_39
timestamp 1644511149
transform 1 0 4692 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_131_51
timestamp 1644511149
transform 1 0 5796 0 -1 73984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_131_55
timestamp 1644511149
transform 1 0 6164 0 -1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_131_57
timestamp 1644511149
transform 1 0 6348 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_131_69
timestamp 1644511149
transform 1 0 7452 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_131_81
timestamp 1644511149
transform 1 0 8556 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_131_93
timestamp 1644511149
transform 1 0 9660 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_131_105
timestamp 1644511149
transform 1 0 10764 0 -1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_131_111
timestamp 1644511149
transform 1 0 11316 0 -1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_131_113
timestamp 1644511149
transform 1 0 11500 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_131_125
timestamp 1644511149
transform 1 0 12604 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_131_137
timestamp 1644511149
transform 1 0 13708 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_131_149
timestamp 1644511149
transform 1 0 14812 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_131_161
timestamp 1644511149
transform 1 0 15916 0 -1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_131_167
timestamp 1644511149
transform 1 0 16468 0 -1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_131_169
timestamp 1644511149
transform 1 0 16652 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_131_181
timestamp 1644511149
transform 1 0 17756 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_131_193
timestamp 1644511149
transform 1 0 18860 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_131_205
timestamp 1644511149
transform 1 0 19964 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_131_217
timestamp 1644511149
transform 1 0 21068 0 -1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_131_223
timestamp 1644511149
transform 1 0 21620 0 -1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_131_225
timestamp 1644511149
transform 1 0 21804 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_131_237
timestamp 1644511149
transform 1 0 22908 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_131_249
timestamp 1644511149
transform 1 0 24012 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_131_261
timestamp 1644511149
transform 1 0 25116 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_131_273
timestamp 1644511149
transform 1 0 26220 0 -1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_131_279
timestamp 1644511149
transform 1 0 26772 0 -1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_131_281
timestamp 1644511149
transform 1 0 26956 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_131_293
timestamp 1644511149
transform 1 0 28060 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_131_305
timestamp 1644511149
transform 1 0 29164 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_131_317
timestamp 1644511149
transform 1 0 30268 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_131_329
timestamp 1644511149
transform 1 0 31372 0 -1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_131_335
timestamp 1644511149
transform 1 0 31924 0 -1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_131_337
timestamp 1644511149
transform 1 0 32108 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_131_349
timestamp 1644511149
transform 1 0 33212 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_131_361
timestamp 1644511149
transform 1 0 34316 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_131_373
timestamp 1644511149
transform 1 0 35420 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_131_385
timestamp 1644511149
transform 1 0 36524 0 -1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_131_391
timestamp 1644511149
transform 1 0 37076 0 -1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_131_393
timestamp 1644511149
transform 1 0 37260 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_131_405
timestamp 1644511149
transform 1 0 38364 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_131_417
timestamp 1644511149
transform 1 0 39468 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_131_429
timestamp 1644511149
transform 1 0 40572 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_131_441
timestamp 1644511149
transform 1 0 41676 0 -1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_131_447
timestamp 1644511149
transform 1 0 42228 0 -1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_131_449
timestamp 1644511149
transform 1 0 42412 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_131_461
timestamp 1644511149
transform 1 0 43516 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_131_473
timestamp 1644511149
transform 1 0 44620 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_131_485
timestamp 1644511149
transform 1 0 45724 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_131_497
timestamp 1644511149
transform 1 0 46828 0 -1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_131_503
timestamp 1644511149
transform 1 0 47380 0 -1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_131_505
timestamp 1644511149
transform 1 0 47564 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_131_517
timestamp 1644511149
transform 1 0 48668 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_131_529
timestamp 1644511149
transform 1 0 49772 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_131_541
timestamp 1644511149
transform 1 0 50876 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_131_553
timestamp 1644511149
transform 1 0 51980 0 -1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_131_559
timestamp 1644511149
transform 1 0 52532 0 -1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_131_561
timestamp 1644511149
transform 1 0 52716 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_131_573
timestamp 1644511149
transform 1 0 53820 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_131_585
timestamp 1644511149
transform 1 0 54924 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_131_597
timestamp 1644511149
transform 1 0 56028 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_131_609
timestamp 1644511149
transform 1 0 57132 0 -1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_131_615
timestamp 1644511149
transform 1 0 57684 0 -1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_131_617
timestamp 1644511149
transform 1 0 57868 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_131_629
timestamp 1644511149
transform 1 0 58972 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_131_641
timestamp 1644511149
transform 1 0 60076 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_131_653
timestamp 1644511149
transform 1 0 61180 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_131_665
timestamp 1644511149
transform 1 0 62284 0 -1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_131_671
timestamp 1644511149
transform 1 0 62836 0 -1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_131_673
timestamp 1644511149
transform 1 0 63020 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_131_685
timestamp 1644511149
transform 1 0 64124 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_131_697
timestamp 1644511149
transform 1 0 65228 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_131_709
timestamp 1644511149
transform 1 0 66332 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_131_721
timestamp 1644511149
transform 1 0 67436 0 -1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_131_727
timestamp 1644511149
transform 1 0 67988 0 -1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_131_729
timestamp 1644511149
transform 1 0 68172 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_131_741
timestamp 1644511149
transform 1 0 69276 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_131_753
timestamp 1644511149
transform 1 0 70380 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_131_765
timestamp 1644511149
transform 1 0 71484 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_131_777
timestamp 1644511149
transform 1 0 72588 0 -1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_131_783
timestamp 1644511149
transform 1 0 73140 0 -1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_131_785
timestamp 1644511149
transform 1 0 73324 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_131_797
timestamp 1644511149
transform 1 0 74428 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_131_809
timestamp 1644511149
transform 1 0 75532 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_131_821
timestamp 1644511149
transform 1 0 76636 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_131_833
timestamp 1644511149
transform 1 0 77740 0 -1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_131_839
timestamp 1644511149
transform 1 0 78292 0 -1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_131_841
timestamp 1644511149
transform 1 0 78476 0 -1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_132_7
timestamp 1644511149
transform 1 0 1748 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_132_19
timestamp 1644511149
transform 1 0 2852 0 1 73984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_132_27
timestamp 1644511149
transform 1 0 3588 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_132_29
timestamp 1644511149
transform 1 0 3772 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_132_41
timestamp 1644511149
transform 1 0 4876 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_132_53
timestamp 1644511149
transform 1 0 5980 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_132_65
timestamp 1644511149
transform 1 0 7084 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_132_77
timestamp 1644511149
transform 1 0 8188 0 1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_132_83
timestamp 1644511149
transform 1 0 8740 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_132_85
timestamp 1644511149
transform 1 0 8924 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_132_97
timestamp 1644511149
transform 1 0 10028 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_132_109
timestamp 1644511149
transform 1 0 11132 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_132_121
timestamp 1644511149
transform 1 0 12236 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_132_133
timestamp 1644511149
transform 1 0 13340 0 1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_132_139
timestamp 1644511149
transform 1 0 13892 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_132_141
timestamp 1644511149
transform 1 0 14076 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_132_153
timestamp 1644511149
transform 1 0 15180 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_132_165
timestamp 1644511149
transform 1 0 16284 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_132_177
timestamp 1644511149
transform 1 0 17388 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_132_189
timestamp 1644511149
transform 1 0 18492 0 1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_132_195
timestamp 1644511149
transform 1 0 19044 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_132_197
timestamp 1644511149
transform 1 0 19228 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_132_209
timestamp 1644511149
transform 1 0 20332 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_132_221
timestamp 1644511149
transform 1 0 21436 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_132_233
timestamp 1644511149
transform 1 0 22540 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_132_245
timestamp 1644511149
transform 1 0 23644 0 1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_132_251
timestamp 1644511149
transform 1 0 24196 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_132_253
timestamp 1644511149
transform 1 0 24380 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_132_265
timestamp 1644511149
transform 1 0 25484 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_132_277
timestamp 1644511149
transform 1 0 26588 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_132_289
timestamp 1644511149
transform 1 0 27692 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_132_301
timestamp 1644511149
transform 1 0 28796 0 1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_132_307
timestamp 1644511149
transform 1 0 29348 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_132_309
timestamp 1644511149
transform 1 0 29532 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_132_321
timestamp 1644511149
transform 1 0 30636 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_132_333
timestamp 1644511149
transform 1 0 31740 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_132_345
timestamp 1644511149
transform 1 0 32844 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_132_357
timestamp 1644511149
transform 1 0 33948 0 1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_132_363
timestamp 1644511149
transform 1 0 34500 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_132_365
timestamp 1644511149
transform 1 0 34684 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_132_377
timestamp 1644511149
transform 1 0 35788 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_132_389
timestamp 1644511149
transform 1 0 36892 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_132_401
timestamp 1644511149
transform 1 0 37996 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_132_413
timestamp 1644511149
transform 1 0 39100 0 1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_132_419
timestamp 1644511149
transform 1 0 39652 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_132_421
timestamp 1644511149
transform 1 0 39836 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_132_433
timestamp 1644511149
transform 1 0 40940 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_132_445
timestamp 1644511149
transform 1 0 42044 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_132_457
timestamp 1644511149
transform 1 0 43148 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_132_469
timestamp 1644511149
transform 1 0 44252 0 1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_132_475
timestamp 1644511149
transform 1 0 44804 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_132_477
timestamp 1644511149
transform 1 0 44988 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_132_489
timestamp 1644511149
transform 1 0 46092 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_132_501
timestamp 1644511149
transform 1 0 47196 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_132_513
timestamp 1644511149
transform 1 0 48300 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_132_525
timestamp 1644511149
transform 1 0 49404 0 1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_132_531
timestamp 1644511149
transform 1 0 49956 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_132_533
timestamp 1644511149
transform 1 0 50140 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_132_545
timestamp 1644511149
transform 1 0 51244 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_132_557
timestamp 1644511149
transform 1 0 52348 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_132_569
timestamp 1644511149
transform 1 0 53452 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_132_581
timestamp 1644511149
transform 1 0 54556 0 1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_132_587
timestamp 1644511149
transform 1 0 55108 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_132_589
timestamp 1644511149
transform 1 0 55292 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_132_601
timestamp 1644511149
transform 1 0 56396 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_132_613
timestamp 1644511149
transform 1 0 57500 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_132_625
timestamp 1644511149
transform 1 0 58604 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_132_637
timestamp 1644511149
transform 1 0 59708 0 1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_132_643
timestamp 1644511149
transform 1 0 60260 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_132_645
timestamp 1644511149
transform 1 0 60444 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_132_657
timestamp 1644511149
transform 1 0 61548 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_132_669
timestamp 1644511149
transform 1 0 62652 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_132_681
timestamp 1644511149
transform 1 0 63756 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_132_693
timestamp 1644511149
transform 1 0 64860 0 1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_132_699
timestamp 1644511149
transform 1 0 65412 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_132_701
timestamp 1644511149
transform 1 0 65596 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_132_713
timestamp 1644511149
transform 1 0 66700 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_132_725
timestamp 1644511149
transform 1 0 67804 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_132_737
timestamp 1644511149
transform 1 0 68908 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_132_749
timestamp 1644511149
transform 1 0 70012 0 1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_132_755
timestamp 1644511149
transform 1 0 70564 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_132_757
timestamp 1644511149
transform 1 0 70748 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_132_769
timestamp 1644511149
transform 1 0 71852 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_132_781
timestamp 1644511149
transform 1 0 72956 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_132_793
timestamp 1644511149
transform 1 0 74060 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_132_805
timestamp 1644511149
transform 1 0 75164 0 1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_132_811
timestamp 1644511149
transform 1 0 75716 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_132_813
timestamp 1644511149
transform 1 0 75900 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_132_825
timestamp 1644511149
transform 1 0 77004 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_132_837
timestamp 1644511149
transform 1 0 78108 0 1 73984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_132_841
timestamp 1644511149
transform 1 0 78476 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_133_3
timestamp 1644511149
transform 1 0 1380 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_133_15
timestamp 1644511149
transform 1 0 2484 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_133_27
timestamp 1644511149
transform 1 0 3588 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_133_39
timestamp 1644511149
transform 1 0 4692 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_133_51
timestamp 1644511149
transform 1 0 5796 0 -1 75072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_133_55
timestamp 1644511149
transform 1 0 6164 0 -1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_133_57
timestamp 1644511149
transform 1 0 6348 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_133_69
timestamp 1644511149
transform 1 0 7452 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_133_81
timestamp 1644511149
transform 1 0 8556 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_133_93
timestamp 1644511149
transform 1 0 9660 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_133_105
timestamp 1644511149
transform 1 0 10764 0 -1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_133_111
timestamp 1644511149
transform 1 0 11316 0 -1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_133_113
timestamp 1644511149
transform 1 0 11500 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_133_125
timestamp 1644511149
transform 1 0 12604 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_133_137
timestamp 1644511149
transform 1 0 13708 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_133_149
timestamp 1644511149
transform 1 0 14812 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_133_161
timestamp 1644511149
transform 1 0 15916 0 -1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_133_167
timestamp 1644511149
transform 1 0 16468 0 -1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_133_169
timestamp 1644511149
transform 1 0 16652 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_133_181
timestamp 1644511149
transform 1 0 17756 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_133_193
timestamp 1644511149
transform 1 0 18860 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_133_205
timestamp 1644511149
transform 1 0 19964 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_133_217
timestamp 1644511149
transform 1 0 21068 0 -1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_133_223
timestamp 1644511149
transform 1 0 21620 0 -1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_133_225
timestamp 1644511149
transform 1 0 21804 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_133_237
timestamp 1644511149
transform 1 0 22908 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_133_249
timestamp 1644511149
transform 1 0 24012 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_133_261
timestamp 1644511149
transform 1 0 25116 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_133_273
timestamp 1644511149
transform 1 0 26220 0 -1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_133_279
timestamp 1644511149
transform 1 0 26772 0 -1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_133_281
timestamp 1644511149
transform 1 0 26956 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_133_293
timestamp 1644511149
transform 1 0 28060 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_133_305
timestamp 1644511149
transform 1 0 29164 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_133_317
timestamp 1644511149
transform 1 0 30268 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_133_329
timestamp 1644511149
transform 1 0 31372 0 -1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_133_335
timestamp 1644511149
transform 1 0 31924 0 -1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_133_337
timestamp 1644511149
transform 1 0 32108 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_133_349
timestamp 1644511149
transform 1 0 33212 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_133_361
timestamp 1644511149
transform 1 0 34316 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_133_373
timestamp 1644511149
transform 1 0 35420 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_133_385
timestamp 1644511149
transform 1 0 36524 0 -1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_133_391
timestamp 1644511149
transform 1 0 37076 0 -1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_133_393
timestamp 1644511149
transform 1 0 37260 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_133_405
timestamp 1644511149
transform 1 0 38364 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_133_417
timestamp 1644511149
transform 1 0 39468 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_133_429
timestamp 1644511149
transform 1 0 40572 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_133_441
timestamp 1644511149
transform 1 0 41676 0 -1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_133_447
timestamp 1644511149
transform 1 0 42228 0 -1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_133_449
timestamp 1644511149
transform 1 0 42412 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_133_461
timestamp 1644511149
transform 1 0 43516 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_133_473
timestamp 1644511149
transform 1 0 44620 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_133_485
timestamp 1644511149
transform 1 0 45724 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_133_497
timestamp 1644511149
transform 1 0 46828 0 -1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_133_503
timestamp 1644511149
transform 1 0 47380 0 -1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_133_505
timestamp 1644511149
transform 1 0 47564 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_133_517
timestamp 1644511149
transform 1 0 48668 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_133_529
timestamp 1644511149
transform 1 0 49772 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_133_541
timestamp 1644511149
transform 1 0 50876 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_133_553
timestamp 1644511149
transform 1 0 51980 0 -1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_133_559
timestamp 1644511149
transform 1 0 52532 0 -1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_133_561
timestamp 1644511149
transform 1 0 52716 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_133_573
timestamp 1644511149
transform 1 0 53820 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_133_585
timestamp 1644511149
transform 1 0 54924 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_133_597
timestamp 1644511149
transform 1 0 56028 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_133_609
timestamp 1644511149
transform 1 0 57132 0 -1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_133_615
timestamp 1644511149
transform 1 0 57684 0 -1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_133_617
timestamp 1644511149
transform 1 0 57868 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_133_629
timestamp 1644511149
transform 1 0 58972 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_133_641
timestamp 1644511149
transform 1 0 60076 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_133_653
timestamp 1644511149
transform 1 0 61180 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_133_665
timestamp 1644511149
transform 1 0 62284 0 -1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_133_671
timestamp 1644511149
transform 1 0 62836 0 -1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_133_673
timestamp 1644511149
transform 1 0 63020 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_133_685
timestamp 1644511149
transform 1 0 64124 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_133_697
timestamp 1644511149
transform 1 0 65228 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_133_709
timestamp 1644511149
transform 1 0 66332 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_133_721
timestamp 1644511149
transform 1 0 67436 0 -1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_133_727
timestamp 1644511149
transform 1 0 67988 0 -1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_133_729
timestamp 1644511149
transform 1 0 68172 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_133_741
timestamp 1644511149
transform 1 0 69276 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_133_753
timestamp 1644511149
transform 1 0 70380 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_133_765
timestamp 1644511149
transform 1 0 71484 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_133_777
timestamp 1644511149
transform 1 0 72588 0 -1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_133_783
timestamp 1644511149
transform 1 0 73140 0 -1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_133_785
timestamp 1644511149
transform 1 0 73324 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_133_797
timestamp 1644511149
transform 1 0 74428 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_133_809
timestamp 1644511149
transform 1 0 75532 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_133_821
timestamp 1644511149
transform 1 0 76636 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_133_833
timestamp 1644511149
transform 1 0 77740 0 -1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_133_839
timestamp 1644511149
transform 1 0 78292 0 -1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_133_841
timestamp 1644511149
transform 1 0 78476 0 -1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_134_3
timestamp 1644511149
transform 1 0 1380 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_134_15
timestamp 1644511149
transform 1 0 2484 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_134_27
timestamp 1644511149
transform 1 0 3588 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_134_29
timestamp 1644511149
transform 1 0 3772 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_134_41
timestamp 1644511149
transform 1 0 4876 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_134_53
timestamp 1644511149
transform 1 0 5980 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_134_65
timestamp 1644511149
transform 1 0 7084 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_134_77
timestamp 1644511149
transform 1 0 8188 0 1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_134_83
timestamp 1644511149
transform 1 0 8740 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_134_85
timestamp 1644511149
transform 1 0 8924 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_134_97
timestamp 1644511149
transform 1 0 10028 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_134_109
timestamp 1644511149
transform 1 0 11132 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_134_121
timestamp 1644511149
transform 1 0 12236 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_134_133
timestamp 1644511149
transform 1 0 13340 0 1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_134_139
timestamp 1644511149
transform 1 0 13892 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_134_141
timestamp 1644511149
transform 1 0 14076 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_134_153
timestamp 1644511149
transform 1 0 15180 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_134_165
timestamp 1644511149
transform 1 0 16284 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_134_177
timestamp 1644511149
transform 1 0 17388 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_134_189
timestamp 1644511149
transform 1 0 18492 0 1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_134_195
timestamp 1644511149
transform 1 0 19044 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_134_197
timestamp 1644511149
transform 1 0 19228 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_134_209
timestamp 1644511149
transform 1 0 20332 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_134_221
timestamp 1644511149
transform 1 0 21436 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_134_233
timestamp 1644511149
transform 1 0 22540 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_134_245
timestamp 1644511149
transform 1 0 23644 0 1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_134_251
timestamp 1644511149
transform 1 0 24196 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_134_253
timestamp 1644511149
transform 1 0 24380 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_134_265
timestamp 1644511149
transform 1 0 25484 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_134_277
timestamp 1644511149
transform 1 0 26588 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_134_289
timestamp 1644511149
transform 1 0 27692 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_134_301
timestamp 1644511149
transform 1 0 28796 0 1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_134_307
timestamp 1644511149
transform 1 0 29348 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_134_309
timestamp 1644511149
transform 1 0 29532 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_134_321
timestamp 1644511149
transform 1 0 30636 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_134_333
timestamp 1644511149
transform 1 0 31740 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_134_345
timestamp 1644511149
transform 1 0 32844 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_134_357
timestamp 1644511149
transform 1 0 33948 0 1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_134_363
timestamp 1644511149
transform 1 0 34500 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_134_365
timestamp 1644511149
transform 1 0 34684 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_134_377
timestamp 1644511149
transform 1 0 35788 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_134_389
timestamp 1644511149
transform 1 0 36892 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_134_401
timestamp 1644511149
transform 1 0 37996 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_134_413
timestamp 1644511149
transform 1 0 39100 0 1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_134_419
timestamp 1644511149
transform 1 0 39652 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_134_421
timestamp 1644511149
transform 1 0 39836 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_134_433
timestamp 1644511149
transform 1 0 40940 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_134_445
timestamp 1644511149
transform 1 0 42044 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_134_457
timestamp 1644511149
transform 1 0 43148 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_134_469
timestamp 1644511149
transform 1 0 44252 0 1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_134_475
timestamp 1644511149
transform 1 0 44804 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_134_477
timestamp 1644511149
transform 1 0 44988 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_134_489
timestamp 1644511149
transform 1 0 46092 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_134_501
timestamp 1644511149
transform 1 0 47196 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_134_513
timestamp 1644511149
transform 1 0 48300 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_134_525
timestamp 1644511149
transform 1 0 49404 0 1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_134_531
timestamp 1644511149
transform 1 0 49956 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_134_533
timestamp 1644511149
transform 1 0 50140 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_134_545
timestamp 1644511149
transform 1 0 51244 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_134_557
timestamp 1644511149
transform 1 0 52348 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_134_569
timestamp 1644511149
transform 1 0 53452 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_134_581
timestamp 1644511149
transform 1 0 54556 0 1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_134_587
timestamp 1644511149
transform 1 0 55108 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_134_589
timestamp 1644511149
transform 1 0 55292 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_134_601
timestamp 1644511149
transform 1 0 56396 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_134_613
timestamp 1644511149
transform 1 0 57500 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_134_625
timestamp 1644511149
transform 1 0 58604 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_134_637
timestamp 1644511149
transform 1 0 59708 0 1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_134_643
timestamp 1644511149
transform 1 0 60260 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_134_645
timestamp 1644511149
transform 1 0 60444 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_134_657
timestamp 1644511149
transform 1 0 61548 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_134_669
timestamp 1644511149
transform 1 0 62652 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_134_681
timestamp 1644511149
transform 1 0 63756 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_134_693
timestamp 1644511149
transform 1 0 64860 0 1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_134_699
timestamp 1644511149
transform 1 0 65412 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_134_701
timestamp 1644511149
transform 1 0 65596 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_134_713
timestamp 1644511149
transform 1 0 66700 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_134_725
timestamp 1644511149
transform 1 0 67804 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_134_737
timestamp 1644511149
transform 1 0 68908 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_134_749
timestamp 1644511149
transform 1 0 70012 0 1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_134_755
timestamp 1644511149
transform 1 0 70564 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_134_757
timestamp 1644511149
transform 1 0 70748 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_134_769
timestamp 1644511149
transform 1 0 71852 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_134_781
timestamp 1644511149
transform 1 0 72956 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_134_793
timestamp 1644511149
transform 1 0 74060 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_134_805
timestamp 1644511149
transform 1 0 75164 0 1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_134_811
timestamp 1644511149
transform 1 0 75716 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_134_813
timestamp 1644511149
transform 1 0 75900 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_134_825
timestamp 1644511149
transform 1 0 77004 0 1 75072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_134_833
timestamp 1644511149
transform 1 0 77740 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_134_838
timestamp 1644511149
transform 1 0 78200 0 1 75072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_135_3
timestamp 1644511149
transform 1 0 1380 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_135_15
timestamp 1644511149
transform 1 0 2484 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_135_27
timestamp 1644511149
transform 1 0 3588 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_135_39
timestamp 1644511149
transform 1 0 4692 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_135_51
timestamp 1644511149
transform 1 0 5796 0 -1 76160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_135_55
timestamp 1644511149
transform 1 0 6164 0 -1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_135_57
timestamp 1644511149
transform 1 0 6348 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_135_69
timestamp 1644511149
transform 1 0 7452 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_135_81
timestamp 1644511149
transform 1 0 8556 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_135_93
timestamp 1644511149
transform 1 0 9660 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_135_105
timestamp 1644511149
transform 1 0 10764 0 -1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_135_111
timestamp 1644511149
transform 1 0 11316 0 -1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_135_113
timestamp 1644511149
transform 1 0 11500 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_135_125
timestamp 1644511149
transform 1 0 12604 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_135_137
timestamp 1644511149
transform 1 0 13708 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_135_149
timestamp 1644511149
transform 1 0 14812 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_135_161
timestamp 1644511149
transform 1 0 15916 0 -1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_135_167
timestamp 1644511149
transform 1 0 16468 0 -1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_135_169
timestamp 1644511149
transform 1 0 16652 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_135_181
timestamp 1644511149
transform 1 0 17756 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_135_193
timestamp 1644511149
transform 1 0 18860 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_135_205
timestamp 1644511149
transform 1 0 19964 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_135_217
timestamp 1644511149
transform 1 0 21068 0 -1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_135_223
timestamp 1644511149
transform 1 0 21620 0 -1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_135_225
timestamp 1644511149
transform 1 0 21804 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_135_237
timestamp 1644511149
transform 1 0 22908 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_135_249
timestamp 1644511149
transform 1 0 24012 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_135_261
timestamp 1644511149
transform 1 0 25116 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_135_273
timestamp 1644511149
transform 1 0 26220 0 -1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_135_279
timestamp 1644511149
transform 1 0 26772 0 -1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_135_281
timestamp 1644511149
transform 1 0 26956 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_135_293
timestamp 1644511149
transform 1 0 28060 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_135_305
timestamp 1644511149
transform 1 0 29164 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_135_317
timestamp 1644511149
transform 1 0 30268 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_135_329
timestamp 1644511149
transform 1 0 31372 0 -1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_135_335
timestamp 1644511149
transform 1 0 31924 0 -1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_135_337
timestamp 1644511149
transform 1 0 32108 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_135_349
timestamp 1644511149
transform 1 0 33212 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_135_361
timestamp 1644511149
transform 1 0 34316 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_135_373
timestamp 1644511149
transform 1 0 35420 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_135_385
timestamp 1644511149
transform 1 0 36524 0 -1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_135_391
timestamp 1644511149
transform 1 0 37076 0 -1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_135_393
timestamp 1644511149
transform 1 0 37260 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_135_405
timestamp 1644511149
transform 1 0 38364 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_135_417
timestamp 1644511149
transform 1 0 39468 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_135_429
timestamp 1644511149
transform 1 0 40572 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_135_441
timestamp 1644511149
transform 1 0 41676 0 -1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_135_447
timestamp 1644511149
transform 1 0 42228 0 -1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_135_449
timestamp 1644511149
transform 1 0 42412 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_135_461
timestamp 1644511149
transform 1 0 43516 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_135_473
timestamp 1644511149
transform 1 0 44620 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_135_485
timestamp 1644511149
transform 1 0 45724 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_135_497
timestamp 1644511149
transform 1 0 46828 0 -1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_135_503
timestamp 1644511149
transform 1 0 47380 0 -1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_135_505
timestamp 1644511149
transform 1 0 47564 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_135_517
timestamp 1644511149
transform 1 0 48668 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_135_529
timestamp 1644511149
transform 1 0 49772 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_135_541
timestamp 1644511149
transform 1 0 50876 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_135_553
timestamp 1644511149
transform 1 0 51980 0 -1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_135_559
timestamp 1644511149
transform 1 0 52532 0 -1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_135_561
timestamp 1644511149
transform 1 0 52716 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_135_573
timestamp 1644511149
transform 1 0 53820 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_135_585
timestamp 1644511149
transform 1 0 54924 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_135_597
timestamp 1644511149
transform 1 0 56028 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_135_609
timestamp 1644511149
transform 1 0 57132 0 -1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_135_615
timestamp 1644511149
transform 1 0 57684 0 -1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_135_617
timestamp 1644511149
transform 1 0 57868 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_135_629
timestamp 1644511149
transform 1 0 58972 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_135_641
timestamp 1644511149
transform 1 0 60076 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_135_653
timestamp 1644511149
transform 1 0 61180 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_135_665
timestamp 1644511149
transform 1 0 62284 0 -1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_135_671
timestamp 1644511149
transform 1 0 62836 0 -1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_135_673
timestamp 1644511149
transform 1 0 63020 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_135_685
timestamp 1644511149
transform 1 0 64124 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_135_697
timestamp 1644511149
transform 1 0 65228 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_135_709
timestamp 1644511149
transform 1 0 66332 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_135_721
timestamp 1644511149
transform 1 0 67436 0 -1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_135_727
timestamp 1644511149
transform 1 0 67988 0 -1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_135_729
timestamp 1644511149
transform 1 0 68172 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_135_741
timestamp 1644511149
transform 1 0 69276 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_135_753
timestamp 1644511149
transform 1 0 70380 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_135_765
timestamp 1644511149
transform 1 0 71484 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_135_777
timestamp 1644511149
transform 1 0 72588 0 -1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_135_783
timestamp 1644511149
transform 1 0 73140 0 -1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_135_785
timestamp 1644511149
transform 1 0 73324 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_135_797
timestamp 1644511149
transform 1 0 74428 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_135_809
timestamp 1644511149
transform 1 0 75532 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_135_821
timestamp 1644511149
transform 1 0 76636 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_135_833
timestamp 1644511149
transform 1 0 77740 0 -1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_135_839
timestamp 1644511149
transform 1 0 78292 0 -1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_135_841
timestamp 1644511149
transform 1 0 78476 0 -1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_136_3
timestamp 1644511149
transform 1 0 1380 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_136_15
timestamp 1644511149
transform 1 0 2484 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_136_27
timestamp 1644511149
transform 1 0 3588 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_136_29
timestamp 1644511149
transform 1 0 3772 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_136_41
timestamp 1644511149
transform 1 0 4876 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_136_53
timestamp 1644511149
transform 1 0 5980 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_136_65
timestamp 1644511149
transform 1 0 7084 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_136_77
timestamp 1644511149
transform 1 0 8188 0 1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_136_83
timestamp 1644511149
transform 1 0 8740 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_136_85
timestamp 1644511149
transform 1 0 8924 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_136_97
timestamp 1644511149
transform 1 0 10028 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_136_109
timestamp 1644511149
transform 1 0 11132 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_136_121
timestamp 1644511149
transform 1 0 12236 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_136_133
timestamp 1644511149
transform 1 0 13340 0 1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_136_139
timestamp 1644511149
transform 1 0 13892 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_136_141
timestamp 1644511149
transform 1 0 14076 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_136_153
timestamp 1644511149
transform 1 0 15180 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_136_165
timestamp 1644511149
transform 1 0 16284 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_136_177
timestamp 1644511149
transform 1 0 17388 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_136_189
timestamp 1644511149
transform 1 0 18492 0 1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_136_195
timestamp 1644511149
transform 1 0 19044 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_136_197
timestamp 1644511149
transform 1 0 19228 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_136_209
timestamp 1644511149
transform 1 0 20332 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_136_221
timestamp 1644511149
transform 1 0 21436 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_136_233
timestamp 1644511149
transform 1 0 22540 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_136_245
timestamp 1644511149
transform 1 0 23644 0 1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_136_251
timestamp 1644511149
transform 1 0 24196 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_136_253
timestamp 1644511149
transform 1 0 24380 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_136_265
timestamp 1644511149
transform 1 0 25484 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_136_277
timestamp 1644511149
transform 1 0 26588 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_136_289
timestamp 1644511149
transform 1 0 27692 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_136_301
timestamp 1644511149
transform 1 0 28796 0 1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_136_307
timestamp 1644511149
transform 1 0 29348 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_136_309
timestamp 1644511149
transform 1 0 29532 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_136_321
timestamp 1644511149
transform 1 0 30636 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_136_333
timestamp 1644511149
transform 1 0 31740 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_136_345
timestamp 1644511149
transform 1 0 32844 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_136_357
timestamp 1644511149
transform 1 0 33948 0 1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_136_363
timestamp 1644511149
transform 1 0 34500 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_136_365
timestamp 1644511149
transform 1 0 34684 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_136_377
timestamp 1644511149
transform 1 0 35788 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_136_389
timestamp 1644511149
transform 1 0 36892 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_136_401
timestamp 1644511149
transform 1 0 37996 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_136_413
timestamp 1644511149
transform 1 0 39100 0 1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_136_419
timestamp 1644511149
transform 1 0 39652 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_136_421
timestamp 1644511149
transform 1 0 39836 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_136_433
timestamp 1644511149
transform 1 0 40940 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_136_445
timestamp 1644511149
transform 1 0 42044 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_136_457
timestamp 1644511149
transform 1 0 43148 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_136_469
timestamp 1644511149
transform 1 0 44252 0 1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_136_475
timestamp 1644511149
transform 1 0 44804 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_136_477
timestamp 1644511149
transform 1 0 44988 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_136_489
timestamp 1644511149
transform 1 0 46092 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_136_501
timestamp 1644511149
transform 1 0 47196 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_136_513
timestamp 1644511149
transform 1 0 48300 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_136_525
timestamp 1644511149
transform 1 0 49404 0 1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_136_531
timestamp 1644511149
transform 1 0 49956 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_136_533
timestamp 1644511149
transform 1 0 50140 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_136_545
timestamp 1644511149
transform 1 0 51244 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_136_557
timestamp 1644511149
transform 1 0 52348 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_136_569
timestamp 1644511149
transform 1 0 53452 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_136_581
timestamp 1644511149
transform 1 0 54556 0 1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_136_587
timestamp 1644511149
transform 1 0 55108 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_136_589
timestamp 1644511149
transform 1 0 55292 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_136_601
timestamp 1644511149
transform 1 0 56396 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_136_613
timestamp 1644511149
transform 1 0 57500 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_136_625
timestamp 1644511149
transform 1 0 58604 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_136_637
timestamp 1644511149
transform 1 0 59708 0 1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_136_643
timestamp 1644511149
transform 1 0 60260 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_136_645
timestamp 1644511149
transform 1 0 60444 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_136_657
timestamp 1644511149
transform 1 0 61548 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_136_669
timestamp 1644511149
transform 1 0 62652 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_136_681
timestamp 1644511149
transform 1 0 63756 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_136_693
timestamp 1644511149
transform 1 0 64860 0 1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_136_699
timestamp 1644511149
transform 1 0 65412 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_136_701
timestamp 1644511149
transform 1 0 65596 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_136_713
timestamp 1644511149
transform 1 0 66700 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_136_725
timestamp 1644511149
transform 1 0 67804 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_136_737
timestamp 1644511149
transform 1 0 68908 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_136_749
timestamp 1644511149
transform 1 0 70012 0 1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_136_755
timestamp 1644511149
transform 1 0 70564 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_136_757
timestamp 1644511149
transform 1 0 70748 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_136_769
timestamp 1644511149
transform 1 0 71852 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_136_781
timestamp 1644511149
transform 1 0 72956 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_136_793
timestamp 1644511149
transform 1 0 74060 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_136_805
timestamp 1644511149
transform 1 0 75164 0 1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_136_811
timestamp 1644511149
transform 1 0 75716 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_136_813
timestamp 1644511149
transform 1 0 75900 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_136_825
timestamp 1644511149
transform 1 0 77004 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_136_837
timestamp 1644511149
transform 1 0 78108 0 1 76160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_136_841
timestamp 1644511149
transform 1 0 78476 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_137_3
timestamp 1644511149
transform 1 0 1380 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_137_15
timestamp 1644511149
transform 1 0 2484 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_137_27
timestamp 1644511149
transform 1 0 3588 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_137_39
timestamp 1644511149
transform 1 0 4692 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_137_51
timestamp 1644511149
transform 1 0 5796 0 -1 77248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_137_55
timestamp 1644511149
transform 1 0 6164 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_137_57
timestamp 1644511149
transform 1 0 6348 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_137_69
timestamp 1644511149
transform 1 0 7452 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_137_81
timestamp 1644511149
transform 1 0 8556 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_137_93
timestamp 1644511149
transform 1 0 9660 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_137_105
timestamp 1644511149
transform 1 0 10764 0 -1 77248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_137_111
timestamp 1644511149
transform 1 0 11316 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_137_113
timestamp 1644511149
transform 1 0 11500 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_137_125
timestamp 1644511149
transform 1 0 12604 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_137_137
timestamp 1644511149
transform 1 0 13708 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_137_149
timestamp 1644511149
transform 1 0 14812 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_137_161
timestamp 1644511149
transform 1 0 15916 0 -1 77248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_137_167
timestamp 1644511149
transform 1 0 16468 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_137_169
timestamp 1644511149
transform 1 0 16652 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_137_181
timestamp 1644511149
transform 1 0 17756 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_137_193
timestamp 1644511149
transform 1 0 18860 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_137_205
timestamp 1644511149
transform 1 0 19964 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_137_217
timestamp 1644511149
transform 1 0 21068 0 -1 77248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_137_223
timestamp 1644511149
transform 1 0 21620 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_137_225
timestamp 1644511149
transform 1 0 21804 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_137_237
timestamp 1644511149
transform 1 0 22908 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_137_249
timestamp 1644511149
transform 1 0 24012 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_137_261
timestamp 1644511149
transform 1 0 25116 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_137_273
timestamp 1644511149
transform 1 0 26220 0 -1 77248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_137_279
timestamp 1644511149
transform 1 0 26772 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_137_281
timestamp 1644511149
transform 1 0 26956 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_137_293
timestamp 1644511149
transform 1 0 28060 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_137_305
timestamp 1644511149
transform 1 0 29164 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_137_317
timestamp 1644511149
transform 1 0 30268 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_137_329
timestamp 1644511149
transform 1 0 31372 0 -1 77248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_137_335
timestamp 1644511149
transform 1 0 31924 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_137_337
timestamp 1644511149
transform 1 0 32108 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_137_349
timestamp 1644511149
transform 1 0 33212 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_137_361
timestamp 1644511149
transform 1 0 34316 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_137_373
timestamp 1644511149
transform 1 0 35420 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_137_385
timestamp 1644511149
transform 1 0 36524 0 -1 77248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_137_391
timestamp 1644511149
transform 1 0 37076 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_137_393
timestamp 1644511149
transform 1 0 37260 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_137_405
timestamp 1644511149
transform 1 0 38364 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_137_417
timestamp 1644511149
transform 1 0 39468 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_137_429
timestamp 1644511149
transform 1 0 40572 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_137_441
timestamp 1644511149
transform 1 0 41676 0 -1 77248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_137_447
timestamp 1644511149
transform 1 0 42228 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_137_449
timestamp 1644511149
transform 1 0 42412 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_137_461
timestamp 1644511149
transform 1 0 43516 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_137_473
timestamp 1644511149
transform 1 0 44620 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_137_485
timestamp 1644511149
transform 1 0 45724 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_137_497
timestamp 1644511149
transform 1 0 46828 0 -1 77248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_137_503
timestamp 1644511149
transform 1 0 47380 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_137_505
timestamp 1644511149
transform 1 0 47564 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_137_517
timestamp 1644511149
transform 1 0 48668 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_137_529
timestamp 1644511149
transform 1 0 49772 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_137_541
timestamp 1644511149
transform 1 0 50876 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_137_553
timestamp 1644511149
transform 1 0 51980 0 -1 77248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_137_559
timestamp 1644511149
transform 1 0 52532 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_137_561
timestamp 1644511149
transform 1 0 52716 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_137_573
timestamp 1644511149
transform 1 0 53820 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_137_585
timestamp 1644511149
transform 1 0 54924 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_137_597
timestamp 1644511149
transform 1 0 56028 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_137_609
timestamp 1644511149
transform 1 0 57132 0 -1 77248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_137_615
timestamp 1644511149
transform 1 0 57684 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_137_617
timestamp 1644511149
transform 1 0 57868 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_137_629
timestamp 1644511149
transform 1 0 58972 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_137_641
timestamp 1644511149
transform 1 0 60076 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_137_653
timestamp 1644511149
transform 1 0 61180 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_137_665
timestamp 1644511149
transform 1 0 62284 0 -1 77248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_137_671
timestamp 1644511149
transform 1 0 62836 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_137_673
timestamp 1644511149
transform 1 0 63020 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_137_685
timestamp 1644511149
transform 1 0 64124 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_137_697
timestamp 1644511149
transform 1 0 65228 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_137_709
timestamp 1644511149
transform 1 0 66332 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_137_721
timestamp 1644511149
transform 1 0 67436 0 -1 77248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_137_727
timestamp 1644511149
transform 1 0 67988 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_137_729
timestamp 1644511149
transform 1 0 68172 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_137_741
timestamp 1644511149
transform 1 0 69276 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_137_753
timestamp 1644511149
transform 1 0 70380 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_137_765
timestamp 1644511149
transform 1 0 71484 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_137_777
timestamp 1644511149
transform 1 0 72588 0 -1 77248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_137_783
timestamp 1644511149
transform 1 0 73140 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_137_785
timestamp 1644511149
transform 1 0 73324 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_137_797
timestamp 1644511149
transform 1 0 74428 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_137_809
timestamp 1644511149
transform 1 0 75532 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_137_821
timestamp 1644511149
transform 1 0 76636 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_137_833
timestamp 1644511149
transform 1 0 77740 0 -1 77248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_137_839
timestamp 1644511149
transform 1 0 78292 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_137_841
timestamp 1644511149
transform 1 0 78476 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_138_3
timestamp 1644511149
transform 1 0 1380 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_138_15
timestamp 1644511149
transform 1 0 2484 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_138_27
timestamp 1644511149
transform 1 0 3588 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_138_29
timestamp 1644511149
transform 1 0 3772 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_138_41
timestamp 1644511149
transform 1 0 4876 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_138_53
timestamp 1644511149
transform 1 0 5980 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_138_65
timestamp 1644511149
transform 1 0 7084 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_138_77
timestamp 1644511149
transform 1 0 8188 0 1 77248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_138_83
timestamp 1644511149
transform 1 0 8740 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_138_85
timestamp 1644511149
transform 1 0 8924 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_138_97
timestamp 1644511149
transform 1 0 10028 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_138_109
timestamp 1644511149
transform 1 0 11132 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_138_121
timestamp 1644511149
transform 1 0 12236 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_138_133
timestamp 1644511149
transform 1 0 13340 0 1 77248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_138_139
timestamp 1644511149
transform 1 0 13892 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_138_141
timestamp 1644511149
transform 1 0 14076 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_138_153
timestamp 1644511149
transform 1 0 15180 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_138_165
timestamp 1644511149
transform 1 0 16284 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_138_177
timestamp 1644511149
transform 1 0 17388 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_138_189
timestamp 1644511149
transform 1 0 18492 0 1 77248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_138_195
timestamp 1644511149
transform 1 0 19044 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_138_197
timestamp 1644511149
transform 1 0 19228 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_138_209
timestamp 1644511149
transform 1 0 20332 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_138_221
timestamp 1644511149
transform 1 0 21436 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_138_233
timestamp 1644511149
transform 1 0 22540 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_138_245
timestamp 1644511149
transform 1 0 23644 0 1 77248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_138_251
timestamp 1644511149
transform 1 0 24196 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_138_253
timestamp 1644511149
transform 1 0 24380 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_138_265
timestamp 1644511149
transform 1 0 25484 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_138_277
timestamp 1644511149
transform 1 0 26588 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_138_289
timestamp 1644511149
transform 1 0 27692 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_138_301
timestamp 1644511149
transform 1 0 28796 0 1 77248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_138_307
timestamp 1644511149
transform 1 0 29348 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_138_309
timestamp 1644511149
transform 1 0 29532 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_138_321
timestamp 1644511149
transform 1 0 30636 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_138_333
timestamp 1644511149
transform 1 0 31740 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_138_345
timestamp 1644511149
transform 1 0 32844 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_138_357
timestamp 1644511149
transform 1 0 33948 0 1 77248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_138_363
timestamp 1644511149
transform 1 0 34500 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_138_365
timestamp 1644511149
transform 1 0 34684 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_138_377
timestamp 1644511149
transform 1 0 35788 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_138_389
timestamp 1644511149
transform 1 0 36892 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_138_401
timestamp 1644511149
transform 1 0 37996 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_138_413
timestamp 1644511149
transform 1 0 39100 0 1 77248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_138_419
timestamp 1644511149
transform 1 0 39652 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_138_421
timestamp 1644511149
transform 1 0 39836 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_138_433
timestamp 1644511149
transform 1 0 40940 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_138_445
timestamp 1644511149
transform 1 0 42044 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_138_457
timestamp 1644511149
transform 1 0 43148 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_138_469
timestamp 1644511149
transform 1 0 44252 0 1 77248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_138_475
timestamp 1644511149
transform 1 0 44804 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_138_477
timestamp 1644511149
transform 1 0 44988 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_138_489
timestamp 1644511149
transform 1 0 46092 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_138_501
timestamp 1644511149
transform 1 0 47196 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_138_513
timestamp 1644511149
transform 1 0 48300 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_138_525
timestamp 1644511149
transform 1 0 49404 0 1 77248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_138_531
timestamp 1644511149
transform 1 0 49956 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_138_533
timestamp 1644511149
transform 1 0 50140 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_138_545
timestamp 1644511149
transform 1 0 51244 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_138_557
timestamp 1644511149
transform 1 0 52348 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_138_569
timestamp 1644511149
transform 1 0 53452 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_138_581
timestamp 1644511149
transform 1 0 54556 0 1 77248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_138_587
timestamp 1644511149
transform 1 0 55108 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_138_589
timestamp 1644511149
transform 1 0 55292 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_138_601
timestamp 1644511149
transform 1 0 56396 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_138_613
timestamp 1644511149
transform 1 0 57500 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_138_625
timestamp 1644511149
transform 1 0 58604 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_138_637
timestamp 1644511149
transform 1 0 59708 0 1 77248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_138_643
timestamp 1644511149
transform 1 0 60260 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_138_645
timestamp 1644511149
transform 1 0 60444 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_138_657
timestamp 1644511149
transform 1 0 61548 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_138_669
timestamp 1644511149
transform 1 0 62652 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_138_681
timestamp 1644511149
transform 1 0 63756 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_138_693
timestamp 1644511149
transform 1 0 64860 0 1 77248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_138_699
timestamp 1644511149
transform 1 0 65412 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_138_701
timestamp 1644511149
transform 1 0 65596 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_138_713
timestamp 1644511149
transform 1 0 66700 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_138_725
timestamp 1644511149
transform 1 0 67804 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_138_737
timestamp 1644511149
transform 1 0 68908 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_138_749
timestamp 1644511149
transform 1 0 70012 0 1 77248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_138_755
timestamp 1644511149
transform 1 0 70564 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_138_757
timestamp 1644511149
transform 1 0 70748 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_138_769
timestamp 1644511149
transform 1 0 71852 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_138_781
timestamp 1644511149
transform 1 0 72956 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_138_793
timestamp 1644511149
transform 1 0 74060 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_138_805
timestamp 1644511149
transform 1 0 75164 0 1 77248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_138_811
timestamp 1644511149
transform 1 0 75716 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_138_813
timestamp 1644511149
transform 1 0 75900 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_138_825
timestamp 1644511149
transform 1 0 77004 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_138_837
timestamp 1644511149
transform 1 0 78108 0 1 77248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_138_841
timestamp 1644511149
transform 1 0 78476 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_139_3
timestamp 1644511149
transform 1 0 1380 0 -1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_139_15
timestamp 1644511149
transform 1 0 2484 0 -1 78336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_139_19
timestamp 1644511149
transform 1 0 2852 0 -1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_139_31
timestamp 1644511149
transform 1 0 3956 0 -1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_139_43
timestamp 1644511149
transform 1 0 5060 0 -1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_139_55
timestamp 1644511149
transform 1 0 6164 0 -1 78336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_139_57
timestamp 1644511149
transform 1 0 6348 0 -1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_139_69
timestamp 1644511149
transform 1 0 7452 0 -1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_139_81
timestamp 1644511149
transform 1 0 8556 0 -1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_139_93
timestamp 1644511149
transform 1 0 9660 0 -1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_139_105
timestamp 1644511149
transform 1 0 10764 0 -1 78336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_139_111
timestamp 1644511149
transform 1 0 11316 0 -1 78336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_139_113
timestamp 1644511149
transform 1 0 11500 0 -1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_139_125
timestamp 1644511149
transform 1 0 12604 0 -1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_139_137
timestamp 1644511149
transform 1 0 13708 0 -1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_139_149
timestamp 1644511149
transform 1 0 14812 0 -1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_139_161
timestamp 1644511149
transform 1 0 15916 0 -1 78336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_139_167
timestamp 1644511149
transform 1 0 16468 0 -1 78336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_139_169
timestamp 1644511149
transform 1 0 16652 0 -1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_139_181
timestamp 1644511149
transform 1 0 17756 0 -1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_139_193
timestamp 1644511149
transform 1 0 18860 0 -1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_139_205
timestamp 1644511149
transform 1 0 19964 0 -1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_139_217
timestamp 1644511149
transform 1 0 21068 0 -1 78336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_139_223
timestamp 1644511149
transform 1 0 21620 0 -1 78336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_139_225
timestamp 1644511149
transform 1 0 21804 0 -1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_139_237
timestamp 1644511149
transform 1 0 22908 0 -1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_139_249
timestamp 1644511149
transform 1 0 24012 0 -1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_139_261
timestamp 1644511149
transform 1 0 25116 0 -1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_139_273
timestamp 1644511149
transform 1 0 26220 0 -1 78336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_139_279
timestamp 1644511149
transform 1 0 26772 0 -1 78336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_139_281
timestamp 1644511149
transform 1 0 26956 0 -1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_139_293
timestamp 1644511149
transform 1 0 28060 0 -1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_139_305
timestamp 1644511149
transform 1 0 29164 0 -1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_139_317
timestamp 1644511149
transform 1 0 30268 0 -1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_139_329
timestamp 1644511149
transform 1 0 31372 0 -1 78336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_139_335
timestamp 1644511149
transform 1 0 31924 0 -1 78336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_139_337
timestamp 1644511149
transform 1 0 32108 0 -1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_139_349
timestamp 1644511149
transform 1 0 33212 0 -1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_139_361
timestamp 1644511149
transform 1 0 34316 0 -1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_139_373
timestamp 1644511149
transform 1 0 35420 0 -1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_139_385
timestamp 1644511149
transform 1 0 36524 0 -1 78336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_139_391
timestamp 1644511149
transform 1 0 37076 0 -1 78336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_139_393
timestamp 1644511149
transform 1 0 37260 0 -1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_139_405
timestamp 1644511149
transform 1 0 38364 0 -1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_139_417
timestamp 1644511149
transform 1 0 39468 0 -1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_139_429
timestamp 1644511149
transform 1 0 40572 0 -1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_139_441
timestamp 1644511149
transform 1 0 41676 0 -1 78336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_139_447
timestamp 1644511149
transform 1 0 42228 0 -1 78336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_139_449
timestamp 1644511149
transform 1 0 42412 0 -1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_139_461
timestamp 1644511149
transform 1 0 43516 0 -1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_139_473
timestamp 1644511149
transform 1 0 44620 0 -1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_139_485
timestamp 1644511149
transform 1 0 45724 0 -1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_139_497
timestamp 1644511149
transform 1 0 46828 0 -1 78336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_139_503
timestamp 1644511149
transform 1 0 47380 0 -1 78336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_139_505
timestamp 1644511149
transform 1 0 47564 0 -1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_139_517
timestamp 1644511149
transform 1 0 48668 0 -1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_139_529
timestamp 1644511149
transform 1 0 49772 0 -1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_139_541
timestamp 1644511149
transform 1 0 50876 0 -1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_139_553
timestamp 1644511149
transform 1 0 51980 0 -1 78336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_139_559
timestamp 1644511149
transform 1 0 52532 0 -1 78336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_139_561
timestamp 1644511149
transform 1 0 52716 0 -1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_139_573
timestamp 1644511149
transform 1 0 53820 0 -1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_139_585
timestamp 1644511149
transform 1 0 54924 0 -1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_139_597
timestamp 1644511149
transform 1 0 56028 0 -1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_139_609
timestamp 1644511149
transform 1 0 57132 0 -1 78336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_139_615
timestamp 1644511149
transform 1 0 57684 0 -1 78336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_139_617
timestamp 1644511149
transform 1 0 57868 0 -1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_139_629
timestamp 1644511149
transform 1 0 58972 0 -1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_139_641
timestamp 1644511149
transform 1 0 60076 0 -1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_139_653
timestamp 1644511149
transform 1 0 61180 0 -1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_139_665
timestamp 1644511149
transform 1 0 62284 0 -1 78336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_139_671
timestamp 1644511149
transform 1 0 62836 0 -1 78336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_139_673
timestamp 1644511149
transform 1 0 63020 0 -1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_139_685
timestamp 1644511149
transform 1 0 64124 0 -1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_139_697
timestamp 1644511149
transform 1 0 65228 0 -1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_139_709
timestamp 1644511149
transform 1 0 66332 0 -1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_139_721
timestamp 1644511149
transform 1 0 67436 0 -1 78336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_139_727
timestamp 1644511149
transform 1 0 67988 0 -1 78336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_139_729
timestamp 1644511149
transform 1 0 68172 0 -1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_139_741
timestamp 1644511149
transform 1 0 69276 0 -1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_139_753
timestamp 1644511149
transform 1 0 70380 0 -1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_139_765
timestamp 1644511149
transform 1 0 71484 0 -1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_139_777
timestamp 1644511149
transform 1 0 72588 0 -1 78336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_139_783
timestamp 1644511149
transform 1 0 73140 0 -1 78336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_139_785
timestamp 1644511149
transform 1 0 73324 0 -1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_139_797
timestamp 1644511149
transform 1 0 74428 0 -1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_139_809
timestamp 1644511149
transform 1 0 75532 0 -1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_139_821
timestamp 1644511149
transform 1 0 76636 0 -1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_139_833
timestamp 1644511149
transform 1 0 77740 0 -1 78336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_139_839
timestamp 1644511149
transform 1 0 78292 0 -1 78336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_139_841
timestamp 1644511149
transform 1 0 78476 0 -1 78336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_140_7
timestamp 1644511149
transform 1 0 1748 0 1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_140_19
timestamp 1644511149
transform 1 0 2852 0 1 78336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_140_27
timestamp 1644511149
transform 1 0 3588 0 1 78336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_140_29
timestamp 1644511149
transform 1 0 3772 0 1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_140_41
timestamp 1644511149
transform 1 0 4876 0 1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_140_53
timestamp 1644511149
transform 1 0 5980 0 1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_140_65
timestamp 1644511149
transform 1 0 7084 0 1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_140_77
timestamp 1644511149
transform 1 0 8188 0 1 78336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_140_83
timestamp 1644511149
transform 1 0 8740 0 1 78336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_140_85
timestamp 1644511149
transform 1 0 8924 0 1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_140_97
timestamp 1644511149
transform 1 0 10028 0 1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_140_109
timestamp 1644511149
transform 1 0 11132 0 1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_140_121
timestamp 1644511149
transform 1 0 12236 0 1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_140_133
timestamp 1644511149
transform 1 0 13340 0 1 78336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_140_139
timestamp 1644511149
transform 1 0 13892 0 1 78336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_140_141
timestamp 1644511149
transform 1 0 14076 0 1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_140_153
timestamp 1644511149
transform 1 0 15180 0 1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_140_165
timestamp 1644511149
transform 1 0 16284 0 1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_140_177
timestamp 1644511149
transform 1 0 17388 0 1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_140_189
timestamp 1644511149
transform 1 0 18492 0 1 78336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_140_195
timestamp 1644511149
transform 1 0 19044 0 1 78336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_140_197
timestamp 1644511149
transform 1 0 19228 0 1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_140_209
timestamp 1644511149
transform 1 0 20332 0 1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_140_221
timestamp 1644511149
transform 1 0 21436 0 1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_140_233
timestamp 1644511149
transform 1 0 22540 0 1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_140_245
timestamp 1644511149
transform 1 0 23644 0 1 78336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_140_251
timestamp 1644511149
transform 1 0 24196 0 1 78336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_140_253
timestamp 1644511149
transform 1 0 24380 0 1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_140_265
timestamp 1644511149
transform 1 0 25484 0 1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_140_277
timestamp 1644511149
transform 1 0 26588 0 1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_140_289
timestamp 1644511149
transform 1 0 27692 0 1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_140_301
timestamp 1644511149
transform 1 0 28796 0 1 78336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_140_307
timestamp 1644511149
transform 1 0 29348 0 1 78336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_140_309
timestamp 1644511149
transform 1 0 29532 0 1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_140_321
timestamp 1644511149
transform 1 0 30636 0 1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_140_333
timestamp 1644511149
transform 1 0 31740 0 1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_140_345
timestamp 1644511149
transform 1 0 32844 0 1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_140_357
timestamp 1644511149
transform 1 0 33948 0 1 78336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_140_363
timestamp 1644511149
transform 1 0 34500 0 1 78336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_140_365
timestamp 1644511149
transform 1 0 34684 0 1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_140_377
timestamp 1644511149
transform 1 0 35788 0 1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_140_389
timestamp 1644511149
transform 1 0 36892 0 1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_140_401
timestamp 1644511149
transform 1 0 37996 0 1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_140_413
timestamp 1644511149
transform 1 0 39100 0 1 78336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_140_419
timestamp 1644511149
transform 1 0 39652 0 1 78336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_140_421
timestamp 1644511149
transform 1 0 39836 0 1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_140_433
timestamp 1644511149
transform 1 0 40940 0 1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_140_445
timestamp 1644511149
transform 1 0 42044 0 1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_140_457
timestamp 1644511149
transform 1 0 43148 0 1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_140_469
timestamp 1644511149
transform 1 0 44252 0 1 78336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_140_475
timestamp 1644511149
transform 1 0 44804 0 1 78336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_140_477
timestamp 1644511149
transform 1 0 44988 0 1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_140_489
timestamp 1644511149
transform 1 0 46092 0 1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_140_501
timestamp 1644511149
transform 1 0 47196 0 1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_140_513
timestamp 1644511149
transform 1 0 48300 0 1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_140_525
timestamp 1644511149
transform 1 0 49404 0 1 78336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_140_531
timestamp 1644511149
transform 1 0 49956 0 1 78336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_140_533
timestamp 1644511149
transform 1 0 50140 0 1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_140_545
timestamp 1644511149
transform 1 0 51244 0 1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_140_557
timestamp 1644511149
transform 1 0 52348 0 1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_140_569
timestamp 1644511149
transform 1 0 53452 0 1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_140_581
timestamp 1644511149
transform 1 0 54556 0 1 78336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_140_587
timestamp 1644511149
transform 1 0 55108 0 1 78336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_140_589
timestamp 1644511149
transform 1 0 55292 0 1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_140_601
timestamp 1644511149
transform 1 0 56396 0 1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_140_613
timestamp 1644511149
transform 1 0 57500 0 1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_140_625
timestamp 1644511149
transform 1 0 58604 0 1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_140_637
timestamp 1644511149
transform 1 0 59708 0 1 78336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_140_643
timestamp 1644511149
transform 1 0 60260 0 1 78336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_140_645
timestamp 1644511149
transform 1 0 60444 0 1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_140_657
timestamp 1644511149
transform 1 0 61548 0 1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_140_669
timestamp 1644511149
transform 1 0 62652 0 1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_140_681
timestamp 1644511149
transform 1 0 63756 0 1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_140_693
timestamp 1644511149
transform 1 0 64860 0 1 78336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_140_699
timestamp 1644511149
transform 1 0 65412 0 1 78336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_140_701
timestamp 1644511149
transform 1 0 65596 0 1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_140_713
timestamp 1644511149
transform 1 0 66700 0 1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_140_725
timestamp 1644511149
transform 1 0 67804 0 1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_140_737
timestamp 1644511149
transform 1 0 68908 0 1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_140_749
timestamp 1644511149
transform 1 0 70012 0 1 78336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_140_755
timestamp 1644511149
transform 1 0 70564 0 1 78336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_140_757
timestamp 1644511149
transform 1 0 70748 0 1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_140_769
timestamp 1644511149
transform 1 0 71852 0 1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_140_781
timestamp 1644511149
transform 1 0 72956 0 1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_140_793
timestamp 1644511149
transform 1 0 74060 0 1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_140_805
timestamp 1644511149
transform 1 0 75164 0 1 78336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_140_811
timestamp 1644511149
transform 1 0 75716 0 1 78336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_140_813
timestamp 1644511149
transform 1 0 75900 0 1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_140_825
timestamp 1644511149
transform 1 0 77004 0 1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_140_837
timestamp 1644511149
transform 1 0 78108 0 1 78336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_140_841
timestamp 1644511149
transform 1 0 78476 0 1 78336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_141_3
timestamp 1644511149
transform 1 0 1380 0 -1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_141_15
timestamp 1644511149
transform 1 0 2484 0 -1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_141_27
timestamp 1644511149
transform 1 0 3588 0 -1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_141_39
timestamp 1644511149
transform 1 0 4692 0 -1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_141_51
timestamp 1644511149
transform 1 0 5796 0 -1 79424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_141_55
timestamp 1644511149
transform 1 0 6164 0 -1 79424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_141_57
timestamp 1644511149
transform 1 0 6348 0 -1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_141_69
timestamp 1644511149
transform 1 0 7452 0 -1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_141_81
timestamp 1644511149
transform 1 0 8556 0 -1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_141_93
timestamp 1644511149
transform 1 0 9660 0 -1 79424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_141_101
timestamp 1644511149
transform 1 0 10396 0 -1 79424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_141_108
timestamp 1644511149
transform 1 0 11040 0 -1 79424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_141_113
timestamp 1644511149
transform 1 0 11500 0 -1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_141_125
timestamp 1644511149
transform 1 0 12604 0 -1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_141_137
timestamp 1644511149
transform 1 0 13708 0 -1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_141_149
timestamp 1644511149
transform 1 0 14812 0 -1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_141_161
timestamp 1644511149
transform 1 0 15916 0 -1 79424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_141_167
timestamp 1644511149
transform 1 0 16468 0 -1 79424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_141_169
timestamp 1644511149
transform 1 0 16652 0 -1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_141_181
timestamp 1644511149
transform 1 0 17756 0 -1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_141_193
timestamp 1644511149
transform 1 0 18860 0 -1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_141_205
timestamp 1644511149
transform 1 0 19964 0 -1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_141_217
timestamp 1644511149
transform 1 0 21068 0 -1 79424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_141_223
timestamp 1644511149
transform 1 0 21620 0 -1 79424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_141_225
timestamp 1644511149
transform 1 0 21804 0 -1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_141_237
timestamp 1644511149
transform 1 0 22908 0 -1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_141_249
timestamp 1644511149
transform 1 0 24012 0 -1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_141_261
timestamp 1644511149
transform 1 0 25116 0 -1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_141_273
timestamp 1644511149
transform 1 0 26220 0 -1 79424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_141_279
timestamp 1644511149
transform 1 0 26772 0 -1 79424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_141_281
timestamp 1644511149
transform 1 0 26956 0 -1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_141_293
timestamp 1644511149
transform 1 0 28060 0 -1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_141_305
timestamp 1644511149
transform 1 0 29164 0 -1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_141_317
timestamp 1644511149
transform 1 0 30268 0 -1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_141_329
timestamp 1644511149
transform 1 0 31372 0 -1 79424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_141_335
timestamp 1644511149
transform 1 0 31924 0 -1 79424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_141_337
timestamp 1644511149
transform 1 0 32108 0 -1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_141_349
timestamp 1644511149
transform 1 0 33212 0 -1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_141_361
timestamp 1644511149
transform 1 0 34316 0 -1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_141_373
timestamp 1644511149
transform 1 0 35420 0 -1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_141_385
timestamp 1644511149
transform 1 0 36524 0 -1 79424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_141_391
timestamp 1644511149
transform 1 0 37076 0 -1 79424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_141_393
timestamp 1644511149
transform 1 0 37260 0 -1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_141_405
timestamp 1644511149
transform 1 0 38364 0 -1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_141_417
timestamp 1644511149
transform 1 0 39468 0 -1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_141_429
timestamp 1644511149
transform 1 0 40572 0 -1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_141_441
timestamp 1644511149
transform 1 0 41676 0 -1 79424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_141_447
timestamp 1644511149
transform 1 0 42228 0 -1 79424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_141_449
timestamp 1644511149
transform 1 0 42412 0 -1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_141_461
timestamp 1644511149
transform 1 0 43516 0 -1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_141_473
timestamp 1644511149
transform 1 0 44620 0 -1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_141_485
timestamp 1644511149
transform 1 0 45724 0 -1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_141_497
timestamp 1644511149
transform 1 0 46828 0 -1 79424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_141_503
timestamp 1644511149
transform 1 0 47380 0 -1 79424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_141_505
timestamp 1644511149
transform 1 0 47564 0 -1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_141_517
timestamp 1644511149
transform 1 0 48668 0 -1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_141_529
timestamp 1644511149
transform 1 0 49772 0 -1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_141_541
timestamp 1644511149
transform 1 0 50876 0 -1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_141_553
timestamp 1644511149
transform 1 0 51980 0 -1 79424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_141_559
timestamp 1644511149
transform 1 0 52532 0 -1 79424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_141_561
timestamp 1644511149
transform 1 0 52716 0 -1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_141_573
timestamp 1644511149
transform 1 0 53820 0 -1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_141_585
timestamp 1644511149
transform 1 0 54924 0 -1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_141_597
timestamp 1644511149
transform 1 0 56028 0 -1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_141_609
timestamp 1644511149
transform 1 0 57132 0 -1 79424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_141_615
timestamp 1644511149
transform 1 0 57684 0 -1 79424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_141_617
timestamp 1644511149
transform 1 0 57868 0 -1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_141_629
timestamp 1644511149
transform 1 0 58972 0 -1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_141_641
timestamp 1644511149
transform 1 0 60076 0 -1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_141_653
timestamp 1644511149
transform 1 0 61180 0 -1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_141_665
timestamp 1644511149
transform 1 0 62284 0 -1 79424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_141_671
timestamp 1644511149
transform 1 0 62836 0 -1 79424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_141_673
timestamp 1644511149
transform 1 0 63020 0 -1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_141_685
timestamp 1644511149
transform 1 0 64124 0 -1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_141_697
timestamp 1644511149
transform 1 0 65228 0 -1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_141_709
timestamp 1644511149
transform 1 0 66332 0 -1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_141_721
timestamp 1644511149
transform 1 0 67436 0 -1 79424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_141_727
timestamp 1644511149
transform 1 0 67988 0 -1 79424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_141_729
timestamp 1644511149
transform 1 0 68172 0 -1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_141_741
timestamp 1644511149
transform 1 0 69276 0 -1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_141_753
timestamp 1644511149
transform 1 0 70380 0 -1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_141_765
timestamp 1644511149
transform 1 0 71484 0 -1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_141_777
timestamp 1644511149
transform 1 0 72588 0 -1 79424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_141_783
timestamp 1644511149
transform 1 0 73140 0 -1 79424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_141_785
timestamp 1644511149
transform 1 0 73324 0 -1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_141_797
timestamp 1644511149
transform 1 0 74428 0 -1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_141_809
timestamp 1644511149
transform 1 0 75532 0 -1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_141_821
timestamp 1644511149
transform 1 0 76636 0 -1 79424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_141_829
timestamp 1644511149
transform 1 0 77372 0 -1 79424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_141_836
timestamp 1644511149
transform 1 0 78016 0 -1 79424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_141_841
timestamp 1644511149
transform 1 0 78476 0 -1 79424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_142_3
timestamp 1644511149
transform 1 0 1380 0 1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_142_15
timestamp 1644511149
transform 1 0 2484 0 1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_142_27
timestamp 1644511149
transform 1 0 3588 0 1 79424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_142_29
timestamp 1644511149
transform 1 0 3772 0 1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_142_41
timestamp 1644511149
transform 1 0 4876 0 1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_142_53
timestamp 1644511149
transform 1 0 5980 0 1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_142_65
timestamp 1644511149
transform 1 0 7084 0 1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_142_77
timestamp 1644511149
transform 1 0 8188 0 1 79424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_142_83
timestamp 1644511149
transform 1 0 8740 0 1 79424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_142_85
timestamp 1644511149
transform 1 0 8924 0 1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_142_97
timestamp 1644511149
transform 1 0 10028 0 1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_142_109
timestamp 1644511149
transform 1 0 11132 0 1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_142_121
timestamp 1644511149
transform 1 0 12236 0 1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_142_133
timestamp 1644511149
transform 1 0 13340 0 1 79424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_142_139
timestamp 1644511149
transform 1 0 13892 0 1 79424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_142_141
timestamp 1644511149
transform 1 0 14076 0 1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_142_153
timestamp 1644511149
transform 1 0 15180 0 1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_142_165
timestamp 1644511149
transform 1 0 16284 0 1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_142_177
timestamp 1644511149
transform 1 0 17388 0 1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_142_189
timestamp 1644511149
transform 1 0 18492 0 1 79424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_142_195
timestamp 1644511149
transform 1 0 19044 0 1 79424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_142_197
timestamp 1644511149
transform 1 0 19228 0 1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_142_209
timestamp 1644511149
transform 1 0 20332 0 1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_142_221
timestamp 1644511149
transform 1 0 21436 0 1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_142_233
timestamp 1644511149
transform 1 0 22540 0 1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_142_245
timestamp 1644511149
transform 1 0 23644 0 1 79424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_142_251
timestamp 1644511149
transform 1 0 24196 0 1 79424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_142_253
timestamp 1644511149
transform 1 0 24380 0 1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_142_265
timestamp 1644511149
transform 1 0 25484 0 1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_142_277
timestamp 1644511149
transform 1 0 26588 0 1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_142_289
timestamp 1644511149
transform 1 0 27692 0 1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_142_301
timestamp 1644511149
transform 1 0 28796 0 1 79424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_142_307
timestamp 1644511149
transform 1 0 29348 0 1 79424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_142_309
timestamp 1644511149
transform 1 0 29532 0 1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_142_321
timestamp 1644511149
transform 1 0 30636 0 1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_142_333
timestamp 1644511149
transform 1 0 31740 0 1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_142_345
timestamp 1644511149
transform 1 0 32844 0 1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_142_357
timestamp 1644511149
transform 1 0 33948 0 1 79424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_142_363
timestamp 1644511149
transform 1 0 34500 0 1 79424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_142_365
timestamp 1644511149
transform 1 0 34684 0 1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_142_377
timestamp 1644511149
transform 1 0 35788 0 1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_142_389
timestamp 1644511149
transform 1 0 36892 0 1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_142_401
timestamp 1644511149
transform 1 0 37996 0 1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_142_413
timestamp 1644511149
transform 1 0 39100 0 1 79424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_142_419
timestamp 1644511149
transform 1 0 39652 0 1 79424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_142_421
timestamp 1644511149
transform 1 0 39836 0 1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_142_433
timestamp 1644511149
transform 1 0 40940 0 1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_142_445
timestamp 1644511149
transform 1 0 42044 0 1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_142_457
timestamp 1644511149
transform 1 0 43148 0 1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_142_469
timestamp 1644511149
transform 1 0 44252 0 1 79424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_142_475
timestamp 1644511149
transform 1 0 44804 0 1 79424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_142_477
timestamp 1644511149
transform 1 0 44988 0 1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_142_489
timestamp 1644511149
transform 1 0 46092 0 1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_142_501
timestamp 1644511149
transform 1 0 47196 0 1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_142_513
timestamp 1644511149
transform 1 0 48300 0 1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_142_525
timestamp 1644511149
transform 1 0 49404 0 1 79424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_142_531
timestamp 1644511149
transform 1 0 49956 0 1 79424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_142_533
timestamp 1644511149
transform 1 0 50140 0 1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_142_545
timestamp 1644511149
transform 1 0 51244 0 1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_142_557
timestamp 1644511149
transform 1 0 52348 0 1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_142_569
timestamp 1644511149
transform 1 0 53452 0 1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_142_581
timestamp 1644511149
transform 1 0 54556 0 1 79424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_142_587
timestamp 1644511149
transform 1 0 55108 0 1 79424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_142_589
timestamp 1644511149
transform 1 0 55292 0 1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_142_601
timestamp 1644511149
transform 1 0 56396 0 1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_142_613
timestamp 1644511149
transform 1 0 57500 0 1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_142_625
timestamp 1644511149
transform 1 0 58604 0 1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_142_637
timestamp 1644511149
transform 1 0 59708 0 1 79424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_142_643
timestamp 1644511149
transform 1 0 60260 0 1 79424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_142_645
timestamp 1644511149
transform 1 0 60444 0 1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_142_657
timestamp 1644511149
transform 1 0 61548 0 1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_142_669
timestamp 1644511149
transform 1 0 62652 0 1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_142_681
timestamp 1644511149
transform 1 0 63756 0 1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_142_693
timestamp 1644511149
transform 1 0 64860 0 1 79424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_142_699
timestamp 1644511149
transform 1 0 65412 0 1 79424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_142_701
timestamp 1644511149
transform 1 0 65596 0 1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_142_713
timestamp 1644511149
transform 1 0 66700 0 1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_142_725
timestamp 1644511149
transform 1 0 67804 0 1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_142_737
timestamp 1644511149
transform 1 0 68908 0 1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_142_749
timestamp 1644511149
transform 1 0 70012 0 1 79424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_142_755
timestamp 1644511149
transform 1 0 70564 0 1 79424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_142_757
timestamp 1644511149
transform 1 0 70748 0 1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_142_769
timestamp 1644511149
transform 1 0 71852 0 1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_142_781
timestamp 1644511149
transform 1 0 72956 0 1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_142_793
timestamp 1644511149
transform 1 0 74060 0 1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_142_805
timestamp 1644511149
transform 1 0 75164 0 1 79424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_142_811
timestamp 1644511149
transform 1 0 75716 0 1 79424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_142_813
timestamp 1644511149
transform 1 0 75900 0 1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_142_825
timestamp 1644511149
transform 1 0 77004 0 1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_142_837
timestamp 1644511149
transform 1 0 78108 0 1 79424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_142_841
timestamp 1644511149
transform 1 0 78476 0 1 79424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_143_3
timestamp 1644511149
transform 1 0 1380 0 -1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_143_15
timestamp 1644511149
transform 1 0 2484 0 -1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_143_27
timestamp 1644511149
transform 1 0 3588 0 -1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_143_39
timestamp 1644511149
transform 1 0 4692 0 -1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_143_51
timestamp 1644511149
transform 1 0 5796 0 -1 80512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_143_55
timestamp 1644511149
transform 1 0 6164 0 -1 80512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_143_57
timestamp 1644511149
transform 1 0 6348 0 -1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_143_69
timestamp 1644511149
transform 1 0 7452 0 -1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_143_81
timestamp 1644511149
transform 1 0 8556 0 -1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_143_93
timestamp 1644511149
transform 1 0 9660 0 -1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_143_105
timestamp 1644511149
transform 1 0 10764 0 -1 80512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_143_111
timestamp 1644511149
transform 1 0 11316 0 -1 80512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_143_113
timestamp 1644511149
transform 1 0 11500 0 -1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_143_125
timestamp 1644511149
transform 1 0 12604 0 -1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_143_137
timestamp 1644511149
transform 1 0 13708 0 -1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_143_149
timestamp 1644511149
transform 1 0 14812 0 -1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_143_161
timestamp 1644511149
transform 1 0 15916 0 -1 80512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_143_167
timestamp 1644511149
transform 1 0 16468 0 -1 80512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_143_169
timestamp 1644511149
transform 1 0 16652 0 -1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_143_181
timestamp 1644511149
transform 1 0 17756 0 -1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_143_193
timestamp 1644511149
transform 1 0 18860 0 -1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_143_205
timestamp 1644511149
transform 1 0 19964 0 -1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_143_217
timestamp 1644511149
transform 1 0 21068 0 -1 80512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_143_223
timestamp 1644511149
transform 1 0 21620 0 -1 80512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_143_225
timestamp 1644511149
transform 1 0 21804 0 -1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_143_237
timestamp 1644511149
transform 1 0 22908 0 -1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_143_249
timestamp 1644511149
transform 1 0 24012 0 -1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_143_261
timestamp 1644511149
transform 1 0 25116 0 -1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_143_273
timestamp 1644511149
transform 1 0 26220 0 -1 80512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_143_279
timestamp 1644511149
transform 1 0 26772 0 -1 80512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_143_281
timestamp 1644511149
transform 1 0 26956 0 -1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_143_293
timestamp 1644511149
transform 1 0 28060 0 -1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_143_305
timestamp 1644511149
transform 1 0 29164 0 -1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_143_317
timestamp 1644511149
transform 1 0 30268 0 -1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_143_329
timestamp 1644511149
transform 1 0 31372 0 -1 80512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_143_335
timestamp 1644511149
transform 1 0 31924 0 -1 80512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_143_337
timestamp 1644511149
transform 1 0 32108 0 -1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_143_349
timestamp 1644511149
transform 1 0 33212 0 -1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_143_361
timestamp 1644511149
transform 1 0 34316 0 -1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_143_373
timestamp 1644511149
transform 1 0 35420 0 -1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_143_385
timestamp 1644511149
transform 1 0 36524 0 -1 80512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_143_391
timestamp 1644511149
transform 1 0 37076 0 -1 80512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_143_393
timestamp 1644511149
transform 1 0 37260 0 -1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_143_405
timestamp 1644511149
transform 1 0 38364 0 -1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_143_417
timestamp 1644511149
transform 1 0 39468 0 -1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_143_429
timestamp 1644511149
transform 1 0 40572 0 -1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_143_441
timestamp 1644511149
transform 1 0 41676 0 -1 80512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_143_447
timestamp 1644511149
transform 1 0 42228 0 -1 80512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_143_449
timestamp 1644511149
transform 1 0 42412 0 -1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_143_461
timestamp 1644511149
transform 1 0 43516 0 -1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_143_473
timestamp 1644511149
transform 1 0 44620 0 -1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_143_485
timestamp 1644511149
transform 1 0 45724 0 -1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_143_497
timestamp 1644511149
transform 1 0 46828 0 -1 80512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_143_503
timestamp 1644511149
transform 1 0 47380 0 -1 80512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_143_505
timestamp 1644511149
transform 1 0 47564 0 -1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_143_517
timestamp 1644511149
transform 1 0 48668 0 -1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_143_529
timestamp 1644511149
transform 1 0 49772 0 -1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_143_541
timestamp 1644511149
transform 1 0 50876 0 -1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_143_553
timestamp 1644511149
transform 1 0 51980 0 -1 80512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_143_559
timestamp 1644511149
transform 1 0 52532 0 -1 80512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_143_561
timestamp 1644511149
transform 1 0 52716 0 -1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_143_573
timestamp 1644511149
transform 1 0 53820 0 -1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_143_585
timestamp 1644511149
transform 1 0 54924 0 -1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_143_597
timestamp 1644511149
transform 1 0 56028 0 -1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_143_609
timestamp 1644511149
transform 1 0 57132 0 -1 80512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_143_615
timestamp 1644511149
transform 1 0 57684 0 -1 80512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_143_617
timestamp 1644511149
transform 1 0 57868 0 -1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_143_629
timestamp 1644511149
transform 1 0 58972 0 -1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_143_641
timestamp 1644511149
transform 1 0 60076 0 -1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_143_653
timestamp 1644511149
transform 1 0 61180 0 -1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_143_665
timestamp 1644511149
transform 1 0 62284 0 -1 80512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_143_671
timestamp 1644511149
transform 1 0 62836 0 -1 80512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_143_673
timestamp 1644511149
transform 1 0 63020 0 -1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_143_685
timestamp 1644511149
transform 1 0 64124 0 -1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_143_697
timestamp 1644511149
transform 1 0 65228 0 -1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_143_709
timestamp 1644511149
transform 1 0 66332 0 -1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_143_721
timestamp 1644511149
transform 1 0 67436 0 -1 80512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_143_727
timestamp 1644511149
transform 1 0 67988 0 -1 80512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_143_729
timestamp 1644511149
transform 1 0 68172 0 -1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_143_741
timestamp 1644511149
transform 1 0 69276 0 -1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_143_753
timestamp 1644511149
transform 1 0 70380 0 -1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_143_765
timestamp 1644511149
transform 1 0 71484 0 -1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_143_777
timestamp 1644511149
transform 1 0 72588 0 -1 80512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_143_783
timestamp 1644511149
transform 1 0 73140 0 -1 80512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_143_785
timestamp 1644511149
transform 1 0 73324 0 -1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_143_797
timestamp 1644511149
transform 1 0 74428 0 -1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_143_809
timestamp 1644511149
transform 1 0 75532 0 -1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_143_821
timestamp 1644511149
transform 1 0 76636 0 -1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_143_833
timestamp 1644511149
transform 1 0 77740 0 -1 80512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_143_839
timestamp 1644511149
transform 1 0 78292 0 -1 80512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_143_841
timestamp 1644511149
transform 1 0 78476 0 -1 80512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_144_3
timestamp 1644511149
transform 1 0 1380 0 1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_144_15
timestamp 1644511149
transform 1 0 2484 0 1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_144_27
timestamp 1644511149
transform 1 0 3588 0 1 80512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_144_29
timestamp 1644511149
transform 1 0 3772 0 1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_144_41
timestamp 1644511149
transform 1 0 4876 0 1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_144_53
timestamp 1644511149
transform 1 0 5980 0 1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_144_65
timestamp 1644511149
transform 1 0 7084 0 1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_144_77
timestamp 1644511149
transform 1 0 8188 0 1 80512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_144_83
timestamp 1644511149
transform 1 0 8740 0 1 80512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_144_85
timestamp 1644511149
transform 1 0 8924 0 1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_144_97
timestamp 1644511149
transform 1 0 10028 0 1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_144_109
timestamp 1644511149
transform 1 0 11132 0 1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_144_121
timestamp 1644511149
transform 1 0 12236 0 1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_144_133
timestamp 1644511149
transform 1 0 13340 0 1 80512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_144_139
timestamp 1644511149
transform 1 0 13892 0 1 80512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_144_141
timestamp 1644511149
transform 1 0 14076 0 1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_144_153
timestamp 1644511149
transform 1 0 15180 0 1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_144_165
timestamp 1644511149
transform 1 0 16284 0 1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_144_177
timestamp 1644511149
transform 1 0 17388 0 1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_144_189
timestamp 1644511149
transform 1 0 18492 0 1 80512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_144_195
timestamp 1644511149
transform 1 0 19044 0 1 80512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_144_197
timestamp 1644511149
transform 1 0 19228 0 1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_144_209
timestamp 1644511149
transform 1 0 20332 0 1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_144_221
timestamp 1644511149
transform 1 0 21436 0 1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_144_233
timestamp 1644511149
transform 1 0 22540 0 1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_144_245
timestamp 1644511149
transform 1 0 23644 0 1 80512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_144_251
timestamp 1644511149
transform 1 0 24196 0 1 80512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_144_253
timestamp 1644511149
transform 1 0 24380 0 1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_144_265
timestamp 1644511149
transform 1 0 25484 0 1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_144_277
timestamp 1644511149
transform 1 0 26588 0 1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_144_289
timestamp 1644511149
transform 1 0 27692 0 1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_144_301
timestamp 1644511149
transform 1 0 28796 0 1 80512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_144_307
timestamp 1644511149
transform 1 0 29348 0 1 80512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_144_309
timestamp 1644511149
transform 1 0 29532 0 1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_144_321
timestamp 1644511149
transform 1 0 30636 0 1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_144_333
timestamp 1644511149
transform 1 0 31740 0 1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_144_345
timestamp 1644511149
transform 1 0 32844 0 1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_144_357
timestamp 1644511149
transform 1 0 33948 0 1 80512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_144_363
timestamp 1644511149
transform 1 0 34500 0 1 80512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_144_365
timestamp 1644511149
transform 1 0 34684 0 1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_144_377
timestamp 1644511149
transform 1 0 35788 0 1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_144_389
timestamp 1644511149
transform 1 0 36892 0 1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_144_401
timestamp 1644511149
transform 1 0 37996 0 1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_144_413
timestamp 1644511149
transform 1 0 39100 0 1 80512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_144_419
timestamp 1644511149
transform 1 0 39652 0 1 80512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_144_421
timestamp 1644511149
transform 1 0 39836 0 1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_144_433
timestamp 1644511149
transform 1 0 40940 0 1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_144_445
timestamp 1644511149
transform 1 0 42044 0 1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_144_457
timestamp 1644511149
transform 1 0 43148 0 1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_144_469
timestamp 1644511149
transform 1 0 44252 0 1 80512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_144_475
timestamp 1644511149
transform 1 0 44804 0 1 80512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_144_477
timestamp 1644511149
transform 1 0 44988 0 1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_144_489
timestamp 1644511149
transform 1 0 46092 0 1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_144_501
timestamp 1644511149
transform 1 0 47196 0 1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_144_513
timestamp 1644511149
transform 1 0 48300 0 1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_144_525
timestamp 1644511149
transform 1 0 49404 0 1 80512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_144_531
timestamp 1644511149
transform 1 0 49956 0 1 80512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_144_533
timestamp 1644511149
transform 1 0 50140 0 1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_144_545
timestamp 1644511149
transform 1 0 51244 0 1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_144_557
timestamp 1644511149
transform 1 0 52348 0 1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_144_569
timestamp 1644511149
transform 1 0 53452 0 1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_144_581
timestamp 1644511149
transform 1 0 54556 0 1 80512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_144_587
timestamp 1644511149
transform 1 0 55108 0 1 80512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_144_589
timestamp 1644511149
transform 1 0 55292 0 1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_144_601
timestamp 1644511149
transform 1 0 56396 0 1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_144_613
timestamp 1644511149
transform 1 0 57500 0 1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_144_625
timestamp 1644511149
transform 1 0 58604 0 1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_144_637
timestamp 1644511149
transform 1 0 59708 0 1 80512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_144_643
timestamp 1644511149
transform 1 0 60260 0 1 80512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_144_645
timestamp 1644511149
transform 1 0 60444 0 1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_144_657
timestamp 1644511149
transform 1 0 61548 0 1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_144_669
timestamp 1644511149
transform 1 0 62652 0 1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_144_681
timestamp 1644511149
transform 1 0 63756 0 1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_144_693
timestamp 1644511149
transform 1 0 64860 0 1 80512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_144_699
timestamp 1644511149
transform 1 0 65412 0 1 80512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_144_701
timestamp 1644511149
transform 1 0 65596 0 1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_144_713
timestamp 1644511149
transform 1 0 66700 0 1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_144_725
timestamp 1644511149
transform 1 0 67804 0 1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_144_737
timestamp 1644511149
transform 1 0 68908 0 1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_144_749
timestamp 1644511149
transform 1 0 70012 0 1 80512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_144_755
timestamp 1644511149
transform 1 0 70564 0 1 80512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_144_757
timestamp 1644511149
transform 1 0 70748 0 1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_144_769
timestamp 1644511149
transform 1 0 71852 0 1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_144_781
timestamp 1644511149
transform 1 0 72956 0 1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_144_793
timestamp 1644511149
transform 1 0 74060 0 1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_144_805
timestamp 1644511149
transform 1 0 75164 0 1 80512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_144_811
timestamp 1644511149
transform 1 0 75716 0 1 80512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_144_813
timestamp 1644511149
transform 1 0 75900 0 1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_144_825
timestamp 1644511149
transform 1 0 77004 0 1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_144_837
timestamp 1644511149
transform 1 0 78108 0 1 80512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_144_841
timestamp 1644511149
transform 1 0 78476 0 1 80512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_145_3
timestamp 1644511149
transform 1 0 1380 0 -1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_145_15
timestamp 1644511149
transform 1 0 2484 0 -1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_145_27
timestamp 1644511149
transform 1 0 3588 0 -1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_145_39
timestamp 1644511149
transform 1 0 4692 0 -1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_145_51
timestamp 1644511149
transform 1 0 5796 0 -1 81600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_145_55
timestamp 1644511149
transform 1 0 6164 0 -1 81600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_145_57
timestamp 1644511149
transform 1 0 6348 0 -1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_145_69
timestamp 1644511149
transform 1 0 7452 0 -1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_145_81
timestamp 1644511149
transform 1 0 8556 0 -1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_145_93
timestamp 1644511149
transform 1 0 9660 0 -1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_145_105
timestamp 1644511149
transform 1 0 10764 0 -1 81600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_145_111
timestamp 1644511149
transform 1 0 11316 0 -1 81600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_145_113
timestamp 1644511149
transform 1 0 11500 0 -1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_145_125
timestamp 1644511149
transform 1 0 12604 0 -1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_145_137
timestamp 1644511149
transform 1 0 13708 0 -1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_145_149
timestamp 1644511149
transform 1 0 14812 0 -1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_145_161
timestamp 1644511149
transform 1 0 15916 0 -1 81600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_145_167
timestamp 1644511149
transform 1 0 16468 0 -1 81600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_145_169
timestamp 1644511149
transform 1 0 16652 0 -1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_145_181
timestamp 1644511149
transform 1 0 17756 0 -1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_145_193
timestamp 1644511149
transform 1 0 18860 0 -1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_145_205
timestamp 1644511149
transform 1 0 19964 0 -1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_145_217
timestamp 1644511149
transform 1 0 21068 0 -1 81600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_145_223
timestamp 1644511149
transform 1 0 21620 0 -1 81600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_145_225
timestamp 1644511149
transform 1 0 21804 0 -1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_145_237
timestamp 1644511149
transform 1 0 22908 0 -1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_145_249
timestamp 1644511149
transform 1 0 24012 0 -1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_145_261
timestamp 1644511149
transform 1 0 25116 0 -1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_145_273
timestamp 1644511149
transform 1 0 26220 0 -1 81600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_145_279
timestamp 1644511149
transform 1 0 26772 0 -1 81600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_145_281
timestamp 1644511149
transform 1 0 26956 0 -1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_145_293
timestamp 1644511149
transform 1 0 28060 0 -1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_145_305
timestamp 1644511149
transform 1 0 29164 0 -1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_145_317
timestamp 1644511149
transform 1 0 30268 0 -1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_145_329
timestamp 1644511149
transform 1 0 31372 0 -1 81600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_145_335
timestamp 1644511149
transform 1 0 31924 0 -1 81600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_145_337
timestamp 1644511149
transform 1 0 32108 0 -1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_145_349
timestamp 1644511149
transform 1 0 33212 0 -1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_145_361
timestamp 1644511149
transform 1 0 34316 0 -1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_145_373
timestamp 1644511149
transform 1 0 35420 0 -1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_145_385
timestamp 1644511149
transform 1 0 36524 0 -1 81600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_145_391
timestamp 1644511149
transform 1 0 37076 0 -1 81600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_145_393
timestamp 1644511149
transform 1 0 37260 0 -1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_145_405
timestamp 1644511149
transform 1 0 38364 0 -1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_145_417
timestamp 1644511149
transform 1 0 39468 0 -1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_145_429
timestamp 1644511149
transform 1 0 40572 0 -1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_145_441
timestamp 1644511149
transform 1 0 41676 0 -1 81600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_145_447
timestamp 1644511149
transform 1 0 42228 0 -1 81600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_145_449
timestamp 1644511149
transform 1 0 42412 0 -1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_145_461
timestamp 1644511149
transform 1 0 43516 0 -1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_145_473
timestamp 1644511149
transform 1 0 44620 0 -1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_145_485
timestamp 1644511149
transform 1 0 45724 0 -1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_145_497
timestamp 1644511149
transform 1 0 46828 0 -1 81600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_145_503
timestamp 1644511149
transform 1 0 47380 0 -1 81600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_145_505
timestamp 1644511149
transform 1 0 47564 0 -1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_145_517
timestamp 1644511149
transform 1 0 48668 0 -1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_145_529
timestamp 1644511149
transform 1 0 49772 0 -1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_145_541
timestamp 1644511149
transform 1 0 50876 0 -1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_145_553
timestamp 1644511149
transform 1 0 51980 0 -1 81600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_145_559
timestamp 1644511149
transform 1 0 52532 0 -1 81600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_145_561
timestamp 1644511149
transform 1 0 52716 0 -1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_145_573
timestamp 1644511149
transform 1 0 53820 0 -1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_145_585
timestamp 1644511149
transform 1 0 54924 0 -1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_145_597
timestamp 1644511149
transform 1 0 56028 0 -1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_145_609
timestamp 1644511149
transform 1 0 57132 0 -1 81600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_145_615
timestamp 1644511149
transform 1 0 57684 0 -1 81600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_145_617
timestamp 1644511149
transform 1 0 57868 0 -1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_145_629
timestamp 1644511149
transform 1 0 58972 0 -1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_145_641
timestamp 1644511149
transform 1 0 60076 0 -1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_145_653
timestamp 1644511149
transform 1 0 61180 0 -1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_145_665
timestamp 1644511149
transform 1 0 62284 0 -1 81600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_145_671
timestamp 1644511149
transform 1 0 62836 0 -1 81600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_145_673
timestamp 1644511149
transform 1 0 63020 0 -1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_145_685
timestamp 1644511149
transform 1 0 64124 0 -1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_145_697
timestamp 1644511149
transform 1 0 65228 0 -1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_145_709
timestamp 1644511149
transform 1 0 66332 0 -1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_145_721
timestamp 1644511149
transform 1 0 67436 0 -1 81600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_145_727
timestamp 1644511149
transform 1 0 67988 0 -1 81600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_145_729
timestamp 1644511149
transform 1 0 68172 0 -1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_145_741
timestamp 1644511149
transform 1 0 69276 0 -1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_145_753
timestamp 1644511149
transform 1 0 70380 0 -1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_145_765
timestamp 1644511149
transform 1 0 71484 0 -1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_145_777
timestamp 1644511149
transform 1 0 72588 0 -1 81600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_145_783
timestamp 1644511149
transform 1 0 73140 0 -1 81600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_145_785
timestamp 1644511149
transform 1 0 73324 0 -1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_145_797
timestamp 1644511149
transform 1 0 74428 0 -1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_145_809
timestamp 1644511149
transform 1 0 75532 0 -1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_145_821
timestamp 1644511149
transform 1 0 76636 0 -1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_145_833
timestamp 1644511149
transform 1 0 77740 0 -1 81600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_145_839
timestamp 1644511149
transform 1 0 78292 0 -1 81600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_145_841
timestamp 1644511149
transform 1 0 78476 0 -1 81600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_146_9
timestamp 1644511149
transform 1 0 1932 0 1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_146_21
timestamp 1644511149
transform 1 0 3036 0 1 81600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_146_27
timestamp 1644511149
transform 1 0 3588 0 1 81600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_146_29
timestamp 1644511149
transform 1 0 3772 0 1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_146_41
timestamp 1644511149
transform 1 0 4876 0 1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_146_53
timestamp 1644511149
transform 1 0 5980 0 1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_146_65
timestamp 1644511149
transform 1 0 7084 0 1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_146_77
timestamp 1644511149
transform 1 0 8188 0 1 81600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_146_83
timestamp 1644511149
transform 1 0 8740 0 1 81600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_146_85
timestamp 1644511149
transform 1 0 8924 0 1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_146_97
timestamp 1644511149
transform 1 0 10028 0 1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_146_109
timestamp 1644511149
transform 1 0 11132 0 1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_146_121
timestamp 1644511149
transform 1 0 12236 0 1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_146_133
timestamp 1644511149
transform 1 0 13340 0 1 81600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_146_139
timestamp 1644511149
transform 1 0 13892 0 1 81600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_146_141
timestamp 1644511149
transform 1 0 14076 0 1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_146_153
timestamp 1644511149
transform 1 0 15180 0 1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_146_165
timestamp 1644511149
transform 1 0 16284 0 1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_146_177
timestamp 1644511149
transform 1 0 17388 0 1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_146_189
timestamp 1644511149
transform 1 0 18492 0 1 81600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_146_195
timestamp 1644511149
transform 1 0 19044 0 1 81600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_146_197
timestamp 1644511149
transform 1 0 19228 0 1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_146_209
timestamp 1644511149
transform 1 0 20332 0 1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_146_221
timestamp 1644511149
transform 1 0 21436 0 1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_146_233
timestamp 1644511149
transform 1 0 22540 0 1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_146_245
timestamp 1644511149
transform 1 0 23644 0 1 81600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_146_251
timestamp 1644511149
transform 1 0 24196 0 1 81600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_146_253
timestamp 1644511149
transform 1 0 24380 0 1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_146_265
timestamp 1644511149
transform 1 0 25484 0 1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_146_277
timestamp 1644511149
transform 1 0 26588 0 1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_146_289
timestamp 1644511149
transform 1 0 27692 0 1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_146_301
timestamp 1644511149
transform 1 0 28796 0 1 81600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_146_307
timestamp 1644511149
transform 1 0 29348 0 1 81600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_146_309
timestamp 1644511149
transform 1 0 29532 0 1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_146_321
timestamp 1644511149
transform 1 0 30636 0 1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_146_333
timestamp 1644511149
transform 1 0 31740 0 1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_146_345
timestamp 1644511149
transform 1 0 32844 0 1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_146_357
timestamp 1644511149
transform 1 0 33948 0 1 81600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_146_363
timestamp 1644511149
transform 1 0 34500 0 1 81600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_146_365
timestamp 1644511149
transform 1 0 34684 0 1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_146_377
timestamp 1644511149
transform 1 0 35788 0 1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_146_389
timestamp 1644511149
transform 1 0 36892 0 1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_146_401
timestamp 1644511149
transform 1 0 37996 0 1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_146_413
timestamp 1644511149
transform 1 0 39100 0 1 81600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_146_419
timestamp 1644511149
transform 1 0 39652 0 1 81600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_146_421
timestamp 1644511149
transform 1 0 39836 0 1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_146_433
timestamp 1644511149
transform 1 0 40940 0 1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_146_445
timestamp 1644511149
transform 1 0 42044 0 1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_146_457
timestamp 1644511149
transform 1 0 43148 0 1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_146_469
timestamp 1644511149
transform 1 0 44252 0 1 81600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_146_475
timestamp 1644511149
transform 1 0 44804 0 1 81600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_146_477
timestamp 1644511149
transform 1 0 44988 0 1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_146_489
timestamp 1644511149
transform 1 0 46092 0 1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_146_501
timestamp 1644511149
transform 1 0 47196 0 1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_146_513
timestamp 1644511149
transform 1 0 48300 0 1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_146_525
timestamp 1644511149
transform 1 0 49404 0 1 81600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_146_531
timestamp 1644511149
transform 1 0 49956 0 1 81600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_146_533
timestamp 1644511149
transform 1 0 50140 0 1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_146_545
timestamp 1644511149
transform 1 0 51244 0 1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_146_557
timestamp 1644511149
transform 1 0 52348 0 1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_146_569
timestamp 1644511149
transform 1 0 53452 0 1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_146_581
timestamp 1644511149
transform 1 0 54556 0 1 81600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_146_587
timestamp 1644511149
transform 1 0 55108 0 1 81600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_146_589
timestamp 1644511149
transform 1 0 55292 0 1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_146_601
timestamp 1644511149
transform 1 0 56396 0 1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_146_613
timestamp 1644511149
transform 1 0 57500 0 1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_146_625
timestamp 1644511149
transform 1 0 58604 0 1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_146_637
timestamp 1644511149
transform 1 0 59708 0 1 81600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_146_643
timestamp 1644511149
transform 1 0 60260 0 1 81600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_146_645
timestamp 1644511149
transform 1 0 60444 0 1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_146_657
timestamp 1644511149
transform 1 0 61548 0 1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_146_669
timestamp 1644511149
transform 1 0 62652 0 1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_146_681
timestamp 1644511149
transform 1 0 63756 0 1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_146_693
timestamp 1644511149
transform 1 0 64860 0 1 81600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_146_699
timestamp 1644511149
transform 1 0 65412 0 1 81600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_146_701
timestamp 1644511149
transform 1 0 65596 0 1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_146_713
timestamp 1644511149
transform 1 0 66700 0 1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_146_725
timestamp 1644511149
transform 1 0 67804 0 1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_146_737
timestamp 1644511149
transform 1 0 68908 0 1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_146_749
timestamp 1644511149
transform 1 0 70012 0 1 81600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_146_755
timestamp 1644511149
transform 1 0 70564 0 1 81600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_146_757
timestamp 1644511149
transform 1 0 70748 0 1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_146_769
timestamp 1644511149
transform 1 0 71852 0 1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_146_781
timestamp 1644511149
transform 1 0 72956 0 1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_146_793
timestamp 1644511149
transform 1 0 74060 0 1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_146_805
timestamp 1644511149
transform 1 0 75164 0 1 81600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_146_811
timestamp 1644511149
transform 1 0 75716 0 1 81600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_146_813
timestamp 1644511149
transform 1 0 75900 0 1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_146_825
timestamp 1644511149
transform 1 0 77004 0 1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_146_837
timestamp 1644511149
transform 1 0 78108 0 1 81600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_146_841
timestamp 1644511149
transform 1 0 78476 0 1 81600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_147_3
timestamp 1644511149
transform 1 0 1380 0 -1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_147_15
timestamp 1644511149
transform 1 0 2484 0 -1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_147_27
timestamp 1644511149
transform 1 0 3588 0 -1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_147_39
timestamp 1644511149
transform 1 0 4692 0 -1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_147_51
timestamp 1644511149
transform 1 0 5796 0 -1 82688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_147_55
timestamp 1644511149
transform 1 0 6164 0 -1 82688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_147_57
timestamp 1644511149
transform 1 0 6348 0 -1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_147_69
timestamp 1644511149
transform 1 0 7452 0 -1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_147_81
timestamp 1644511149
transform 1 0 8556 0 -1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_147_93
timestamp 1644511149
transform 1 0 9660 0 -1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_147_105
timestamp 1644511149
transform 1 0 10764 0 -1 82688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_147_111
timestamp 1644511149
transform 1 0 11316 0 -1 82688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_147_113
timestamp 1644511149
transform 1 0 11500 0 -1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_147_125
timestamp 1644511149
transform 1 0 12604 0 -1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_147_137
timestamp 1644511149
transform 1 0 13708 0 -1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_147_149
timestamp 1644511149
transform 1 0 14812 0 -1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_147_161
timestamp 1644511149
transform 1 0 15916 0 -1 82688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_147_167
timestamp 1644511149
transform 1 0 16468 0 -1 82688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_147_169
timestamp 1644511149
transform 1 0 16652 0 -1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_147_181
timestamp 1644511149
transform 1 0 17756 0 -1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_147_193
timestamp 1644511149
transform 1 0 18860 0 -1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_147_205
timestamp 1644511149
transform 1 0 19964 0 -1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_147_217
timestamp 1644511149
transform 1 0 21068 0 -1 82688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_147_223
timestamp 1644511149
transform 1 0 21620 0 -1 82688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_147_225
timestamp 1644511149
transform 1 0 21804 0 -1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_147_237
timestamp 1644511149
transform 1 0 22908 0 -1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_147_249
timestamp 1644511149
transform 1 0 24012 0 -1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_147_261
timestamp 1644511149
transform 1 0 25116 0 -1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_147_273
timestamp 1644511149
transform 1 0 26220 0 -1 82688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_147_279
timestamp 1644511149
transform 1 0 26772 0 -1 82688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_147_281
timestamp 1644511149
transform 1 0 26956 0 -1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_147_293
timestamp 1644511149
transform 1 0 28060 0 -1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_147_305
timestamp 1644511149
transform 1 0 29164 0 -1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_147_317
timestamp 1644511149
transform 1 0 30268 0 -1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_147_329
timestamp 1644511149
transform 1 0 31372 0 -1 82688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_147_335
timestamp 1644511149
transform 1 0 31924 0 -1 82688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_147_337
timestamp 1644511149
transform 1 0 32108 0 -1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_147_349
timestamp 1644511149
transform 1 0 33212 0 -1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_147_361
timestamp 1644511149
transform 1 0 34316 0 -1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_147_373
timestamp 1644511149
transform 1 0 35420 0 -1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_147_385
timestamp 1644511149
transform 1 0 36524 0 -1 82688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_147_391
timestamp 1644511149
transform 1 0 37076 0 -1 82688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_147_393
timestamp 1644511149
transform 1 0 37260 0 -1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_147_405
timestamp 1644511149
transform 1 0 38364 0 -1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_147_417
timestamp 1644511149
transform 1 0 39468 0 -1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_147_429
timestamp 1644511149
transform 1 0 40572 0 -1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_147_441
timestamp 1644511149
transform 1 0 41676 0 -1 82688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_147_447
timestamp 1644511149
transform 1 0 42228 0 -1 82688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_147_449
timestamp 1644511149
transform 1 0 42412 0 -1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_147_461
timestamp 1644511149
transform 1 0 43516 0 -1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_147_473
timestamp 1644511149
transform 1 0 44620 0 -1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_147_485
timestamp 1644511149
transform 1 0 45724 0 -1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_147_497
timestamp 1644511149
transform 1 0 46828 0 -1 82688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_147_503
timestamp 1644511149
transform 1 0 47380 0 -1 82688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_147_505
timestamp 1644511149
transform 1 0 47564 0 -1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_147_517
timestamp 1644511149
transform 1 0 48668 0 -1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_147_529
timestamp 1644511149
transform 1 0 49772 0 -1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_147_541
timestamp 1644511149
transform 1 0 50876 0 -1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_147_553
timestamp 1644511149
transform 1 0 51980 0 -1 82688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_147_559
timestamp 1644511149
transform 1 0 52532 0 -1 82688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_147_561
timestamp 1644511149
transform 1 0 52716 0 -1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_147_573
timestamp 1644511149
transform 1 0 53820 0 -1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_147_585
timestamp 1644511149
transform 1 0 54924 0 -1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_147_597
timestamp 1644511149
transform 1 0 56028 0 -1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_147_609
timestamp 1644511149
transform 1 0 57132 0 -1 82688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_147_615
timestamp 1644511149
transform 1 0 57684 0 -1 82688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_147_617
timestamp 1644511149
transform 1 0 57868 0 -1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_147_629
timestamp 1644511149
transform 1 0 58972 0 -1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_147_641
timestamp 1644511149
transform 1 0 60076 0 -1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_147_653
timestamp 1644511149
transform 1 0 61180 0 -1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_147_665
timestamp 1644511149
transform 1 0 62284 0 -1 82688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_147_671
timestamp 1644511149
transform 1 0 62836 0 -1 82688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_147_673
timestamp 1644511149
transform 1 0 63020 0 -1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_147_685
timestamp 1644511149
transform 1 0 64124 0 -1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_147_697
timestamp 1644511149
transform 1 0 65228 0 -1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_147_709
timestamp 1644511149
transform 1 0 66332 0 -1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_147_721
timestamp 1644511149
transform 1 0 67436 0 -1 82688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_147_727
timestamp 1644511149
transform 1 0 67988 0 -1 82688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_147_729
timestamp 1644511149
transform 1 0 68172 0 -1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_147_741
timestamp 1644511149
transform 1 0 69276 0 -1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_147_753
timestamp 1644511149
transform 1 0 70380 0 -1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_147_765
timestamp 1644511149
transform 1 0 71484 0 -1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_147_777
timestamp 1644511149
transform 1 0 72588 0 -1 82688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_147_783
timestamp 1644511149
transform 1 0 73140 0 -1 82688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_147_785
timestamp 1644511149
transform 1 0 73324 0 -1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_147_797
timestamp 1644511149
transform 1 0 74428 0 -1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_147_809
timestamp 1644511149
transform 1 0 75532 0 -1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_147_821
timestamp 1644511149
transform 1 0 76636 0 -1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_147_833
timestamp 1644511149
transform 1 0 77740 0 -1 82688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_147_839
timestamp 1644511149
transform 1 0 78292 0 -1 82688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_147_841
timestamp 1644511149
transform 1 0 78476 0 -1 82688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_148_3
timestamp 1644511149
transform 1 0 1380 0 1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_148_15
timestamp 1644511149
transform 1 0 2484 0 1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_148_27
timestamp 1644511149
transform 1 0 3588 0 1 82688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_148_29
timestamp 1644511149
transform 1 0 3772 0 1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_148_41
timestamp 1644511149
transform 1 0 4876 0 1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_148_53
timestamp 1644511149
transform 1 0 5980 0 1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_148_65
timestamp 1644511149
transform 1 0 7084 0 1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_148_77
timestamp 1644511149
transform 1 0 8188 0 1 82688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_148_83
timestamp 1644511149
transform 1 0 8740 0 1 82688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_148_85
timestamp 1644511149
transform 1 0 8924 0 1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_148_97
timestamp 1644511149
transform 1 0 10028 0 1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_148_109
timestamp 1644511149
transform 1 0 11132 0 1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_148_121
timestamp 1644511149
transform 1 0 12236 0 1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_148_133
timestamp 1644511149
transform 1 0 13340 0 1 82688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_148_139
timestamp 1644511149
transform 1 0 13892 0 1 82688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_148_141
timestamp 1644511149
transform 1 0 14076 0 1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_148_153
timestamp 1644511149
transform 1 0 15180 0 1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_148_165
timestamp 1644511149
transform 1 0 16284 0 1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_148_177
timestamp 1644511149
transform 1 0 17388 0 1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_148_189
timestamp 1644511149
transform 1 0 18492 0 1 82688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_148_195
timestamp 1644511149
transform 1 0 19044 0 1 82688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_148_197
timestamp 1644511149
transform 1 0 19228 0 1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_148_209
timestamp 1644511149
transform 1 0 20332 0 1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_148_221
timestamp 1644511149
transform 1 0 21436 0 1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_148_233
timestamp 1644511149
transform 1 0 22540 0 1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_148_245
timestamp 1644511149
transform 1 0 23644 0 1 82688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_148_251
timestamp 1644511149
transform 1 0 24196 0 1 82688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_148_253
timestamp 1644511149
transform 1 0 24380 0 1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_148_265
timestamp 1644511149
transform 1 0 25484 0 1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_148_277
timestamp 1644511149
transform 1 0 26588 0 1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_148_289
timestamp 1644511149
transform 1 0 27692 0 1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_148_301
timestamp 1644511149
transform 1 0 28796 0 1 82688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_148_307
timestamp 1644511149
transform 1 0 29348 0 1 82688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_148_309
timestamp 1644511149
transform 1 0 29532 0 1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_148_321
timestamp 1644511149
transform 1 0 30636 0 1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_148_333
timestamp 1644511149
transform 1 0 31740 0 1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_148_345
timestamp 1644511149
transform 1 0 32844 0 1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_148_357
timestamp 1644511149
transform 1 0 33948 0 1 82688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_148_363
timestamp 1644511149
transform 1 0 34500 0 1 82688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_148_365
timestamp 1644511149
transform 1 0 34684 0 1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_148_377
timestamp 1644511149
transform 1 0 35788 0 1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_148_389
timestamp 1644511149
transform 1 0 36892 0 1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_148_401
timestamp 1644511149
transform 1 0 37996 0 1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_148_413
timestamp 1644511149
transform 1 0 39100 0 1 82688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_148_419
timestamp 1644511149
transform 1 0 39652 0 1 82688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_148_421
timestamp 1644511149
transform 1 0 39836 0 1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_148_433
timestamp 1644511149
transform 1 0 40940 0 1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_148_445
timestamp 1644511149
transform 1 0 42044 0 1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_148_457
timestamp 1644511149
transform 1 0 43148 0 1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_148_469
timestamp 1644511149
transform 1 0 44252 0 1 82688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_148_475
timestamp 1644511149
transform 1 0 44804 0 1 82688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_148_477
timestamp 1644511149
transform 1 0 44988 0 1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_148_489
timestamp 1644511149
transform 1 0 46092 0 1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_148_501
timestamp 1644511149
transform 1 0 47196 0 1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_148_513
timestamp 1644511149
transform 1 0 48300 0 1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_148_525
timestamp 1644511149
transform 1 0 49404 0 1 82688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_148_531
timestamp 1644511149
transform 1 0 49956 0 1 82688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_148_533
timestamp 1644511149
transform 1 0 50140 0 1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_148_545
timestamp 1644511149
transform 1 0 51244 0 1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_148_557
timestamp 1644511149
transform 1 0 52348 0 1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_148_569
timestamp 1644511149
transform 1 0 53452 0 1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_148_581
timestamp 1644511149
transform 1 0 54556 0 1 82688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_148_587
timestamp 1644511149
transform 1 0 55108 0 1 82688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_148_589
timestamp 1644511149
transform 1 0 55292 0 1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_148_601
timestamp 1644511149
transform 1 0 56396 0 1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_148_613
timestamp 1644511149
transform 1 0 57500 0 1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_148_625
timestamp 1644511149
transform 1 0 58604 0 1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_148_637
timestamp 1644511149
transform 1 0 59708 0 1 82688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_148_643
timestamp 1644511149
transform 1 0 60260 0 1 82688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_148_645
timestamp 1644511149
transform 1 0 60444 0 1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_148_657
timestamp 1644511149
transform 1 0 61548 0 1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_148_669
timestamp 1644511149
transform 1 0 62652 0 1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_148_681
timestamp 1644511149
transform 1 0 63756 0 1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_148_693
timestamp 1644511149
transform 1 0 64860 0 1 82688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_148_699
timestamp 1644511149
transform 1 0 65412 0 1 82688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_148_701
timestamp 1644511149
transform 1 0 65596 0 1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_148_713
timestamp 1644511149
transform 1 0 66700 0 1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_148_725
timestamp 1644511149
transform 1 0 67804 0 1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_148_737
timestamp 1644511149
transform 1 0 68908 0 1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_148_749
timestamp 1644511149
transform 1 0 70012 0 1 82688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_148_755
timestamp 1644511149
transform 1 0 70564 0 1 82688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_148_757
timestamp 1644511149
transform 1 0 70748 0 1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_148_769
timestamp 1644511149
transform 1 0 71852 0 1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_148_781
timestamp 1644511149
transform 1 0 72956 0 1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_148_793
timestamp 1644511149
transform 1 0 74060 0 1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_148_805
timestamp 1644511149
transform 1 0 75164 0 1 82688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_148_811
timestamp 1644511149
transform 1 0 75716 0 1 82688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_148_813
timestamp 1644511149
transform 1 0 75900 0 1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_148_825
timestamp 1644511149
transform 1 0 77004 0 1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_148_837
timestamp 1644511149
transform 1 0 78108 0 1 82688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_148_841
timestamp 1644511149
transform 1 0 78476 0 1 82688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_149_3
timestamp 1644511149
transform 1 0 1380 0 -1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_149_15
timestamp 1644511149
transform 1 0 2484 0 -1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_149_27
timestamp 1644511149
transform 1 0 3588 0 -1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_149_39
timestamp 1644511149
transform 1 0 4692 0 -1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_149_51
timestamp 1644511149
transform 1 0 5796 0 -1 83776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_149_55
timestamp 1644511149
transform 1 0 6164 0 -1 83776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_149_57
timestamp 1644511149
transform 1 0 6348 0 -1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_149_69
timestamp 1644511149
transform 1 0 7452 0 -1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_149_81
timestamp 1644511149
transform 1 0 8556 0 -1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_149_93
timestamp 1644511149
transform 1 0 9660 0 -1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_149_105
timestamp 1644511149
transform 1 0 10764 0 -1 83776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_149_111
timestamp 1644511149
transform 1 0 11316 0 -1 83776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_149_113
timestamp 1644511149
transform 1 0 11500 0 -1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_149_125
timestamp 1644511149
transform 1 0 12604 0 -1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_149_137
timestamp 1644511149
transform 1 0 13708 0 -1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_149_149
timestamp 1644511149
transform 1 0 14812 0 -1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_149_161
timestamp 1644511149
transform 1 0 15916 0 -1 83776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_149_167
timestamp 1644511149
transform 1 0 16468 0 -1 83776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_149_169
timestamp 1644511149
transform 1 0 16652 0 -1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_149_181
timestamp 1644511149
transform 1 0 17756 0 -1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_149_193
timestamp 1644511149
transform 1 0 18860 0 -1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_149_205
timestamp 1644511149
transform 1 0 19964 0 -1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_149_217
timestamp 1644511149
transform 1 0 21068 0 -1 83776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_149_223
timestamp 1644511149
transform 1 0 21620 0 -1 83776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_149_225
timestamp 1644511149
transform 1 0 21804 0 -1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_149_237
timestamp 1644511149
transform 1 0 22908 0 -1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_149_249
timestamp 1644511149
transform 1 0 24012 0 -1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_149_261
timestamp 1644511149
transform 1 0 25116 0 -1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_149_273
timestamp 1644511149
transform 1 0 26220 0 -1 83776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_149_279
timestamp 1644511149
transform 1 0 26772 0 -1 83776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_149_281
timestamp 1644511149
transform 1 0 26956 0 -1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_149_293
timestamp 1644511149
transform 1 0 28060 0 -1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_149_305
timestamp 1644511149
transform 1 0 29164 0 -1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_149_317
timestamp 1644511149
transform 1 0 30268 0 -1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_149_329
timestamp 1644511149
transform 1 0 31372 0 -1 83776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_149_335
timestamp 1644511149
transform 1 0 31924 0 -1 83776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_149_337
timestamp 1644511149
transform 1 0 32108 0 -1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_149_349
timestamp 1644511149
transform 1 0 33212 0 -1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_149_361
timestamp 1644511149
transform 1 0 34316 0 -1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_149_373
timestamp 1644511149
transform 1 0 35420 0 -1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_149_385
timestamp 1644511149
transform 1 0 36524 0 -1 83776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_149_391
timestamp 1644511149
transform 1 0 37076 0 -1 83776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_149_393
timestamp 1644511149
transform 1 0 37260 0 -1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_149_405
timestamp 1644511149
transform 1 0 38364 0 -1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_149_417
timestamp 1644511149
transform 1 0 39468 0 -1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_149_429
timestamp 1644511149
transform 1 0 40572 0 -1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_149_441
timestamp 1644511149
transform 1 0 41676 0 -1 83776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_149_447
timestamp 1644511149
transform 1 0 42228 0 -1 83776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_149_449
timestamp 1644511149
transform 1 0 42412 0 -1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_149_461
timestamp 1644511149
transform 1 0 43516 0 -1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_149_473
timestamp 1644511149
transform 1 0 44620 0 -1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_149_485
timestamp 1644511149
transform 1 0 45724 0 -1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_149_497
timestamp 1644511149
transform 1 0 46828 0 -1 83776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_149_503
timestamp 1644511149
transform 1 0 47380 0 -1 83776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_149_505
timestamp 1644511149
transform 1 0 47564 0 -1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_149_517
timestamp 1644511149
transform 1 0 48668 0 -1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_149_529
timestamp 1644511149
transform 1 0 49772 0 -1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_149_541
timestamp 1644511149
transform 1 0 50876 0 -1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_149_553
timestamp 1644511149
transform 1 0 51980 0 -1 83776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_149_559
timestamp 1644511149
transform 1 0 52532 0 -1 83776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_149_561
timestamp 1644511149
transform 1 0 52716 0 -1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_149_573
timestamp 1644511149
transform 1 0 53820 0 -1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_149_585
timestamp 1644511149
transform 1 0 54924 0 -1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_149_597
timestamp 1644511149
transform 1 0 56028 0 -1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_149_609
timestamp 1644511149
transform 1 0 57132 0 -1 83776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_149_615
timestamp 1644511149
transform 1 0 57684 0 -1 83776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_149_617
timestamp 1644511149
transform 1 0 57868 0 -1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_149_629
timestamp 1644511149
transform 1 0 58972 0 -1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_149_641
timestamp 1644511149
transform 1 0 60076 0 -1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_149_653
timestamp 1644511149
transform 1 0 61180 0 -1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_149_665
timestamp 1644511149
transform 1 0 62284 0 -1 83776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_149_671
timestamp 1644511149
transform 1 0 62836 0 -1 83776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_149_673
timestamp 1644511149
transform 1 0 63020 0 -1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_149_685
timestamp 1644511149
transform 1 0 64124 0 -1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_149_697
timestamp 1644511149
transform 1 0 65228 0 -1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_149_709
timestamp 1644511149
transform 1 0 66332 0 -1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_149_721
timestamp 1644511149
transform 1 0 67436 0 -1 83776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_149_727
timestamp 1644511149
transform 1 0 67988 0 -1 83776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_149_729
timestamp 1644511149
transform 1 0 68172 0 -1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_149_741
timestamp 1644511149
transform 1 0 69276 0 -1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_149_753
timestamp 1644511149
transform 1 0 70380 0 -1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_149_765
timestamp 1644511149
transform 1 0 71484 0 -1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_149_777
timestamp 1644511149
transform 1 0 72588 0 -1 83776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_149_783
timestamp 1644511149
transform 1 0 73140 0 -1 83776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_149_785
timestamp 1644511149
transform 1 0 73324 0 -1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_149_797
timestamp 1644511149
transform 1 0 74428 0 -1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_149_809
timestamp 1644511149
transform 1 0 75532 0 -1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_149_821
timestamp 1644511149
transform 1 0 76636 0 -1 83776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_149_829
timestamp 1644511149
transform 1 0 77372 0 -1 83776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_149_836
timestamp 1644511149
transform 1 0 78016 0 -1 83776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_149_841
timestamp 1644511149
transform 1 0 78476 0 -1 83776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_150_3
timestamp 1644511149
transform 1 0 1380 0 1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_150_15
timestamp 1644511149
transform 1 0 2484 0 1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_150_27
timestamp 1644511149
transform 1 0 3588 0 1 83776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_150_29
timestamp 1644511149
transform 1 0 3772 0 1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_150_41
timestamp 1644511149
transform 1 0 4876 0 1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_150_53
timestamp 1644511149
transform 1 0 5980 0 1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_150_65
timestamp 1644511149
transform 1 0 7084 0 1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_150_77
timestamp 1644511149
transform 1 0 8188 0 1 83776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_150_83
timestamp 1644511149
transform 1 0 8740 0 1 83776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_150_85
timestamp 1644511149
transform 1 0 8924 0 1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_150_97
timestamp 1644511149
transform 1 0 10028 0 1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_150_109
timestamp 1644511149
transform 1 0 11132 0 1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_150_121
timestamp 1644511149
transform 1 0 12236 0 1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_150_133
timestamp 1644511149
transform 1 0 13340 0 1 83776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_150_139
timestamp 1644511149
transform 1 0 13892 0 1 83776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_150_141
timestamp 1644511149
transform 1 0 14076 0 1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_150_153
timestamp 1644511149
transform 1 0 15180 0 1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_150_165
timestamp 1644511149
transform 1 0 16284 0 1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_150_177
timestamp 1644511149
transform 1 0 17388 0 1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_150_189
timestamp 1644511149
transform 1 0 18492 0 1 83776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_150_195
timestamp 1644511149
transform 1 0 19044 0 1 83776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_150_197
timestamp 1644511149
transform 1 0 19228 0 1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_150_209
timestamp 1644511149
transform 1 0 20332 0 1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_150_221
timestamp 1644511149
transform 1 0 21436 0 1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_150_233
timestamp 1644511149
transform 1 0 22540 0 1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_150_245
timestamp 1644511149
transform 1 0 23644 0 1 83776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_150_251
timestamp 1644511149
transform 1 0 24196 0 1 83776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_150_253
timestamp 1644511149
transform 1 0 24380 0 1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_150_265
timestamp 1644511149
transform 1 0 25484 0 1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_150_277
timestamp 1644511149
transform 1 0 26588 0 1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_150_289
timestamp 1644511149
transform 1 0 27692 0 1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_150_301
timestamp 1644511149
transform 1 0 28796 0 1 83776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_150_307
timestamp 1644511149
transform 1 0 29348 0 1 83776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_150_309
timestamp 1644511149
transform 1 0 29532 0 1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_150_321
timestamp 1644511149
transform 1 0 30636 0 1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_150_333
timestamp 1644511149
transform 1 0 31740 0 1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_150_345
timestamp 1644511149
transform 1 0 32844 0 1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_150_357
timestamp 1644511149
transform 1 0 33948 0 1 83776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_150_363
timestamp 1644511149
transform 1 0 34500 0 1 83776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_150_365
timestamp 1644511149
transform 1 0 34684 0 1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_150_377
timestamp 1644511149
transform 1 0 35788 0 1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_150_389
timestamp 1644511149
transform 1 0 36892 0 1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_150_401
timestamp 1644511149
transform 1 0 37996 0 1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_150_413
timestamp 1644511149
transform 1 0 39100 0 1 83776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_150_419
timestamp 1644511149
transform 1 0 39652 0 1 83776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_150_421
timestamp 1644511149
transform 1 0 39836 0 1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_150_433
timestamp 1644511149
transform 1 0 40940 0 1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_150_445
timestamp 1644511149
transform 1 0 42044 0 1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_150_457
timestamp 1644511149
transform 1 0 43148 0 1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_150_469
timestamp 1644511149
transform 1 0 44252 0 1 83776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_150_475
timestamp 1644511149
transform 1 0 44804 0 1 83776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_150_477
timestamp 1644511149
transform 1 0 44988 0 1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_150_489
timestamp 1644511149
transform 1 0 46092 0 1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_150_501
timestamp 1644511149
transform 1 0 47196 0 1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_150_513
timestamp 1644511149
transform 1 0 48300 0 1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_150_525
timestamp 1644511149
transform 1 0 49404 0 1 83776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_150_531
timestamp 1644511149
transform 1 0 49956 0 1 83776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_150_533
timestamp 1644511149
transform 1 0 50140 0 1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_150_545
timestamp 1644511149
transform 1 0 51244 0 1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_150_557
timestamp 1644511149
transform 1 0 52348 0 1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_150_569
timestamp 1644511149
transform 1 0 53452 0 1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_150_581
timestamp 1644511149
transform 1 0 54556 0 1 83776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_150_587
timestamp 1644511149
transform 1 0 55108 0 1 83776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_150_589
timestamp 1644511149
transform 1 0 55292 0 1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_150_601
timestamp 1644511149
transform 1 0 56396 0 1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_150_613
timestamp 1644511149
transform 1 0 57500 0 1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_150_625
timestamp 1644511149
transform 1 0 58604 0 1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_150_637
timestamp 1644511149
transform 1 0 59708 0 1 83776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_150_643
timestamp 1644511149
transform 1 0 60260 0 1 83776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_150_645
timestamp 1644511149
transform 1 0 60444 0 1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_150_657
timestamp 1644511149
transform 1 0 61548 0 1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_150_669
timestamp 1644511149
transform 1 0 62652 0 1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_150_681
timestamp 1644511149
transform 1 0 63756 0 1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_150_693
timestamp 1644511149
transform 1 0 64860 0 1 83776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_150_699
timestamp 1644511149
transform 1 0 65412 0 1 83776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_150_701
timestamp 1644511149
transform 1 0 65596 0 1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_150_713
timestamp 1644511149
transform 1 0 66700 0 1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_150_725
timestamp 1644511149
transform 1 0 67804 0 1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_150_737
timestamp 1644511149
transform 1 0 68908 0 1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_150_749
timestamp 1644511149
transform 1 0 70012 0 1 83776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_150_755
timestamp 1644511149
transform 1 0 70564 0 1 83776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_150_757
timestamp 1644511149
transform 1 0 70748 0 1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_150_769
timestamp 1644511149
transform 1 0 71852 0 1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_150_781
timestamp 1644511149
transform 1 0 72956 0 1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_150_793
timestamp 1644511149
transform 1 0 74060 0 1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_150_805
timestamp 1644511149
transform 1 0 75164 0 1 83776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_150_811
timestamp 1644511149
transform 1 0 75716 0 1 83776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_150_813
timestamp 1644511149
transform 1 0 75900 0 1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_150_825
timestamp 1644511149
transform 1 0 77004 0 1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_150_837
timestamp 1644511149
transform 1 0 78108 0 1 83776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_150_841
timestamp 1644511149
transform 1 0 78476 0 1 83776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_151_3
timestamp 1644511149
transform 1 0 1380 0 -1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_151_15
timestamp 1644511149
transform 1 0 2484 0 -1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_151_27
timestamp 1644511149
transform 1 0 3588 0 -1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_151_39
timestamp 1644511149
transform 1 0 4692 0 -1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_151_51
timestamp 1644511149
transform 1 0 5796 0 -1 84864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_151_55
timestamp 1644511149
transform 1 0 6164 0 -1 84864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_151_57
timestamp 1644511149
transform 1 0 6348 0 -1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_151_69
timestamp 1644511149
transform 1 0 7452 0 -1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_151_81
timestamp 1644511149
transform 1 0 8556 0 -1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_151_93
timestamp 1644511149
transform 1 0 9660 0 -1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_151_105
timestamp 1644511149
transform 1 0 10764 0 -1 84864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_151_111
timestamp 1644511149
transform 1 0 11316 0 -1 84864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_151_113
timestamp 1644511149
transform 1 0 11500 0 -1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_151_125
timestamp 1644511149
transform 1 0 12604 0 -1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_151_137
timestamp 1644511149
transform 1 0 13708 0 -1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_151_149
timestamp 1644511149
transform 1 0 14812 0 -1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_151_161
timestamp 1644511149
transform 1 0 15916 0 -1 84864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_151_167
timestamp 1644511149
transform 1 0 16468 0 -1 84864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_151_169
timestamp 1644511149
transform 1 0 16652 0 -1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_151_181
timestamp 1644511149
transform 1 0 17756 0 -1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_151_193
timestamp 1644511149
transform 1 0 18860 0 -1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_151_205
timestamp 1644511149
transform 1 0 19964 0 -1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_151_217
timestamp 1644511149
transform 1 0 21068 0 -1 84864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_151_223
timestamp 1644511149
transform 1 0 21620 0 -1 84864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_151_225
timestamp 1644511149
transform 1 0 21804 0 -1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_151_237
timestamp 1644511149
transform 1 0 22908 0 -1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_151_249
timestamp 1644511149
transform 1 0 24012 0 -1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_151_261
timestamp 1644511149
transform 1 0 25116 0 -1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_151_273
timestamp 1644511149
transform 1 0 26220 0 -1 84864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_151_279
timestamp 1644511149
transform 1 0 26772 0 -1 84864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_151_281
timestamp 1644511149
transform 1 0 26956 0 -1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_151_293
timestamp 1644511149
transform 1 0 28060 0 -1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_151_305
timestamp 1644511149
transform 1 0 29164 0 -1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_151_317
timestamp 1644511149
transform 1 0 30268 0 -1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_151_329
timestamp 1644511149
transform 1 0 31372 0 -1 84864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_151_335
timestamp 1644511149
transform 1 0 31924 0 -1 84864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_151_337
timestamp 1644511149
transform 1 0 32108 0 -1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_151_349
timestamp 1644511149
transform 1 0 33212 0 -1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_151_361
timestamp 1644511149
transform 1 0 34316 0 -1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_151_373
timestamp 1644511149
transform 1 0 35420 0 -1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_151_385
timestamp 1644511149
transform 1 0 36524 0 -1 84864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_151_391
timestamp 1644511149
transform 1 0 37076 0 -1 84864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_151_393
timestamp 1644511149
transform 1 0 37260 0 -1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_151_405
timestamp 1644511149
transform 1 0 38364 0 -1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_151_417
timestamp 1644511149
transform 1 0 39468 0 -1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_151_429
timestamp 1644511149
transform 1 0 40572 0 -1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_151_441
timestamp 1644511149
transform 1 0 41676 0 -1 84864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_151_447
timestamp 1644511149
transform 1 0 42228 0 -1 84864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_151_449
timestamp 1644511149
transform 1 0 42412 0 -1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_151_461
timestamp 1644511149
transform 1 0 43516 0 -1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_151_473
timestamp 1644511149
transform 1 0 44620 0 -1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_151_485
timestamp 1644511149
transform 1 0 45724 0 -1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_151_497
timestamp 1644511149
transform 1 0 46828 0 -1 84864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_151_503
timestamp 1644511149
transform 1 0 47380 0 -1 84864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_151_505
timestamp 1644511149
transform 1 0 47564 0 -1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_151_517
timestamp 1644511149
transform 1 0 48668 0 -1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_151_529
timestamp 1644511149
transform 1 0 49772 0 -1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_151_541
timestamp 1644511149
transform 1 0 50876 0 -1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_151_553
timestamp 1644511149
transform 1 0 51980 0 -1 84864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_151_559
timestamp 1644511149
transform 1 0 52532 0 -1 84864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_151_561
timestamp 1644511149
transform 1 0 52716 0 -1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_151_573
timestamp 1644511149
transform 1 0 53820 0 -1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_151_585
timestamp 1644511149
transform 1 0 54924 0 -1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_151_597
timestamp 1644511149
transform 1 0 56028 0 -1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_151_609
timestamp 1644511149
transform 1 0 57132 0 -1 84864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_151_615
timestamp 1644511149
transform 1 0 57684 0 -1 84864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_151_617
timestamp 1644511149
transform 1 0 57868 0 -1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_151_629
timestamp 1644511149
transform 1 0 58972 0 -1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_151_641
timestamp 1644511149
transform 1 0 60076 0 -1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_151_653
timestamp 1644511149
transform 1 0 61180 0 -1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_151_665
timestamp 1644511149
transform 1 0 62284 0 -1 84864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_151_671
timestamp 1644511149
transform 1 0 62836 0 -1 84864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_151_673
timestamp 1644511149
transform 1 0 63020 0 -1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_151_685
timestamp 1644511149
transform 1 0 64124 0 -1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_151_697
timestamp 1644511149
transform 1 0 65228 0 -1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_151_709
timestamp 1644511149
transform 1 0 66332 0 -1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_151_721
timestamp 1644511149
transform 1 0 67436 0 -1 84864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_151_727
timestamp 1644511149
transform 1 0 67988 0 -1 84864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_151_729
timestamp 1644511149
transform 1 0 68172 0 -1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_151_741
timestamp 1644511149
transform 1 0 69276 0 -1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_151_753
timestamp 1644511149
transform 1 0 70380 0 -1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_151_765
timestamp 1644511149
transform 1 0 71484 0 -1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_151_777
timestamp 1644511149
transform 1 0 72588 0 -1 84864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_151_783
timestamp 1644511149
transform 1 0 73140 0 -1 84864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_151_785
timestamp 1644511149
transform 1 0 73324 0 -1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_151_797
timestamp 1644511149
transform 1 0 74428 0 -1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_151_809
timestamp 1644511149
transform 1 0 75532 0 -1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_151_821
timestamp 1644511149
transform 1 0 76636 0 -1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_151_833
timestamp 1644511149
transform 1 0 77740 0 -1 84864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_151_839
timestamp 1644511149
transform 1 0 78292 0 -1 84864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_151_841
timestamp 1644511149
transform 1 0 78476 0 -1 84864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_152_3
timestamp 1644511149
transform 1 0 1380 0 1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_152_15
timestamp 1644511149
transform 1 0 2484 0 1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_152_27
timestamp 1644511149
transform 1 0 3588 0 1 84864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_152_29
timestamp 1644511149
transform 1 0 3772 0 1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_152_41
timestamp 1644511149
transform 1 0 4876 0 1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_152_53
timestamp 1644511149
transform 1 0 5980 0 1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_152_65
timestamp 1644511149
transform 1 0 7084 0 1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_152_77
timestamp 1644511149
transform 1 0 8188 0 1 84864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_152_83
timestamp 1644511149
transform 1 0 8740 0 1 84864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_152_85
timestamp 1644511149
transform 1 0 8924 0 1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_152_97
timestamp 1644511149
transform 1 0 10028 0 1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_152_109
timestamp 1644511149
transform 1 0 11132 0 1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_152_121
timestamp 1644511149
transform 1 0 12236 0 1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_152_133
timestamp 1644511149
transform 1 0 13340 0 1 84864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_152_139
timestamp 1644511149
transform 1 0 13892 0 1 84864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_152_141
timestamp 1644511149
transform 1 0 14076 0 1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_152_153
timestamp 1644511149
transform 1 0 15180 0 1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_152_165
timestamp 1644511149
transform 1 0 16284 0 1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_152_177
timestamp 1644511149
transform 1 0 17388 0 1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_152_189
timestamp 1644511149
transform 1 0 18492 0 1 84864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_152_195
timestamp 1644511149
transform 1 0 19044 0 1 84864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_152_197
timestamp 1644511149
transform 1 0 19228 0 1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_152_209
timestamp 1644511149
transform 1 0 20332 0 1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_152_221
timestamp 1644511149
transform 1 0 21436 0 1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_152_233
timestamp 1644511149
transform 1 0 22540 0 1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_152_245
timestamp 1644511149
transform 1 0 23644 0 1 84864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_152_251
timestamp 1644511149
transform 1 0 24196 0 1 84864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_152_253
timestamp 1644511149
transform 1 0 24380 0 1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_152_265
timestamp 1644511149
transform 1 0 25484 0 1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_152_277
timestamp 1644511149
transform 1 0 26588 0 1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_152_289
timestamp 1644511149
transform 1 0 27692 0 1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_152_301
timestamp 1644511149
transform 1 0 28796 0 1 84864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_152_307
timestamp 1644511149
transform 1 0 29348 0 1 84864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_152_309
timestamp 1644511149
transform 1 0 29532 0 1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_152_321
timestamp 1644511149
transform 1 0 30636 0 1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_152_333
timestamp 1644511149
transform 1 0 31740 0 1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_152_345
timestamp 1644511149
transform 1 0 32844 0 1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_152_357
timestamp 1644511149
transform 1 0 33948 0 1 84864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_152_363
timestamp 1644511149
transform 1 0 34500 0 1 84864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_152_365
timestamp 1644511149
transform 1 0 34684 0 1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_152_377
timestamp 1644511149
transform 1 0 35788 0 1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_152_389
timestamp 1644511149
transform 1 0 36892 0 1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_152_401
timestamp 1644511149
transform 1 0 37996 0 1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_152_413
timestamp 1644511149
transform 1 0 39100 0 1 84864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_152_419
timestamp 1644511149
transform 1 0 39652 0 1 84864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_152_421
timestamp 1644511149
transform 1 0 39836 0 1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_152_433
timestamp 1644511149
transform 1 0 40940 0 1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_152_445
timestamp 1644511149
transform 1 0 42044 0 1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_152_457
timestamp 1644511149
transform 1 0 43148 0 1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_152_469
timestamp 1644511149
transform 1 0 44252 0 1 84864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_152_475
timestamp 1644511149
transform 1 0 44804 0 1 84864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_152_477
timestamp 1644511149
transform 1 0 44988 0 1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_152_489
timestamp 1644511149
transform 1 0 46092 0 1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_152_501
timestamp 1644511149
transform 1 0 47196 0 1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_152_513
timestamp 1644511149
transform 1 0 48300 0 1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_152_525
timestamp 1644511149
transform 1 0 49404 0 1 84864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_152_531
timestamp 1644511149
transform 1 0 49956 0 1 84864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_152_533
timestamp 1644511149
transform 1 0 50140 0 1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_152_545
timestamp 1644511149
transform 1 0 51244 0 1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_152_557
timestamp 1644511149
transform 1 0 52348 0 1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_152_569
timestamp 1644511149
transform 1 0 53452 0 1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_152_581
timestamp 1644511149
transform 1 0 54556 0 1 84864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_152_587
timestamp 1644511149
transform 1 0 55108 0 1 84864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_152_589
timestamp 1644511149
transform 1 0 55292 0 1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_152_601
timestamp 1644511149
transform 1 0 56396 0 1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_152_613
timestamp 1644511149
transform 1 0 57500 0 1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_152_625
timestamp 1644511149
transform 1 0 58604 0 1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_152_637
timestamp 1644511149
transform 1 0 59708 0 1 84864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_152_643
timestamp 1644511149
transform 1 0 60260 0 1 84864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_152_645
timestamp 1644511149
transform 1 0 60444 0 1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_152_657
timestamp 1644511149
transform 1 0 61548 0 1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_152_669
timestamp 1644511149
transform 1 0 62652 0 1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_152_681
timestamp 1644511149
transform 1 0 63756 0 1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_152_693
timestamp 1644511149
transform 1 0 64860 0 1 84864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_152_699
timestamp 1644511149
transform 1 0 65412 0 1 84864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_152_701
timestamp 1644511149
transform 1 0 65596 0 1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_152_713
timestamp 1644511149
transform 1 0 66700 0 1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_152_725
timestamp 1644511149
transform 1 0 67804 0 1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_152_737
timestamp 1644511149
transform 1 0 68908 0 1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_152_749
timestamp 1644511149
transform 1 0 70012 0 1 84864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_152_755
timestamp 1644511149
transform 1 0 70564 0 1 84864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_152_757
timestamp 1644511149
transform 1 0 70748 0 1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_152_769
timestamp 1644511149
transform 1 0 71852 0 1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_152_781
timestamp 1644511149
transform 1 0 72956 0 1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_152_793
timestamp 1644511149
transform 1 0 74060 0 1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_152_805
timestamp 1644511149
transform 1 0 75164 0 1 84864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_152_811
timestamp 1644511149
transform 1 0 75716 0 1 84864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_152_813
timestamp 1644511149
transform 1 0 75900 0 1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_152_825
timestamp 1644511149
transform 1 0 77004 0 1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_152_837
timestamp 1644511149
transform 1 0 78108 0 1 84864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_152_841
timestamp 1644511149
transform 1 0 78476 0 1 84864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_153_3
timestamp 1644511149
transform 1 0 1380 0 -1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_153_15
timestamp 1644511149
transform 1 0 2484 0 -1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_153_27
timestamp 1644511149
transform 1 0 3588 0 -1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_153_39
timestamp 1644511149
transform 1 0 4692 0 -1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_153_51
timestamp 1644511149
transform 1 0 5796 0 -1 85952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_153_55
timestamp 1644511149
transform 1 0 6164 0 -1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_153_57
timestamp 1644511149
transform 1 0 6348 0 -1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_153_69
timestamp 1644511149
transform 1 0 7452 0 -1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_153_81
timestamp 1644511149
transform 1 0 8556 0 -1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_153_93
timestamp 1644511149
transform 1 0 9660 0 -1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_153_105
timestamp 1644511149
transform 1 0 10764 0 -1 85952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_153_111
timestamp 1644511149
transform 1 0 11316 0 -1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_153_113
timestamp 1644511149
transform 1 0 11500 0 -1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_153_125
timestamp 1644511149
transform 1 0 12604 0 -1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_153_137
timestamp 1644511149
transform 1 0 13708 0 -1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_153_149
timestamp 1644511149
transform 1 0 14812 0 -1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_153_161
timestamp 1644511149
transform 1 0 15916 0 -1 85952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_153_167
timestamp 1644511149
transform 1 0 16468 0 -1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_153_169
timestamp 1644511149
transform 1 0 16652 0 -1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_153_181
timestamp 1644511149
transform 1 0 17756 0 -1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_153_193
timestamp 1644511149
transform 1 0 18860 0 -1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_153_205
timestamp 1644511149
transform 1 0 19964 0 -1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_153_217
timestamp 1644511149
transform 1 0 21068 0 -1 85952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_153_223
timestamp 1644511149
transform 1 0 21620 0 -1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_153_225
timestamp 1644511149
transform 1 0 21804 0 -1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_153_237
timestamp 1644511149
transform 1 0 22908 0 -1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_153_249
timestamp 1644511149
transform 1 0 24012 0 -1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_153_261
timestamp 1644511149
transform 1 0 25116 0 -1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_153_273
timestamp 1644511149
transform 1 0 26220 0 -1 85952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_153_279
timestamp 1644511149
transform 1 0 26772 0 -1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_153_281
timestamp 1644511149
transform 1 0 26956 0 -1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_153_293
timestamp 1644511149
transform 1 0 28060 0 -1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_153_305
timestamp 1644511149
transform 1 0 29164 0 -1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_153_317
timestamp 1644511149
transform 1 0 30268 0 -1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_153_329
timestamp 1644511149
transform 1 0 31372 0 -1 85952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_153_335
timestamp 1644511149
transform 1 0 31924 0 -1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_153_337
timestamp 1644511149
transform 1 0 32108 0 -1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_153_349
timestamp 1644511149
transform 1 0 33212 0 -1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_153_361
timestamp 1644511149
transform 1 0 34316 0 -1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_153_373
timestamp 1644511149
transform 1 0 35420 0 -1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_153_385
timestamp 1644511149
transform 1 0 36524 0 -1 85952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_153_391
timestamp 1644511149
transform 1 0 37076 0 -1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_153_393
timestamp 1644511149
transform 1 0 37260 0 -1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_153_405
timestamp 1644511149
transform 1 0 38364 0 -1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_153_417
timestamp 1644511149
transform 1 0 39468 0 -1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_153_429
timestamp 1644511149
transform 1 0 40572 0 -1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_153_441
timestamp 1644511149
transform 1 0 41676 0 -1 85952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_153_447
timestamp 1644511149
transform 1 0 42228 0 -1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_153_449
timestamp 1644511149
transform 1 0 42412 0 -1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_153_461
timestamp 1644511149
transform 1 0 43516 0 -1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_153_473
timestamp 1644511149
transform 1 0 44620 0 -1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_153_485
timestamp 1644511149
transform 1 0 45724 0 -1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_153_497
timestamp 1644511149
transform 1 0 46828 0 -1 85952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_153_503
timestamp 1644511149
transform 1 0 47380 0 -1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_153_505
timestamp 1644511149
transform 1 0 47564 0 -1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_153_517
timestamp 1644511149
transform 1 0 48668 0 -1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_153_529
timestamp 1644511149
transform 1 0 49772 0 -1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_153_541
timestamp 1644511149
transform 1 0 50876 0 -1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_153_553
timestamp 1644511149
transform 1 0 51980 0 -1 85952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_153_559
timestamp 1644511149
transform 1 0 52532 0 -1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_153_561
timestamp 1644511149
transform 1 0 52716 0 -1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_153_573
timestamp 1644511149
transform 1 0 53820 0 -1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_153_585
timestamp 1644511149
transform 1 0 54924 0 -1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_153_597
timestamp 1644511149
transform 1 0 56028 0 -1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_153_609
timestamp 1644511149
transform 1 0 57132 0 -1 85952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_153_615
timestamp 1644511149
transform 1 0 57684 0 -1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_153_617
timestamp 1644511149
transform 1 0 57868 0 -1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_153_629
timestamp 1644511149
transform 1 0 58972 0 -1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_153_641
timestamp 1644511149
transform 1 0 60076 0 -1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_153_653
timestamp 1644511149
transform 1 0 61180 0 -1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_153_665
timestamp 1644511149
transform 1 0 62284 0 -1 85952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_153_671
timestamp 1644511149
transform 1 0 62836 0 -1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_153_673
timestamp 1644511149
transform 1 0 63020 0 -1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_153_685
timestamp 1644511149
transform 1 0 64124 0 -1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_153_697
timestamp 1644511149
transform 1 0 65228 0 -1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_153_709
timestamp 1644511149
transform 1 0 66332 0 -1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_153_721
timestamp 1644511149
transform 1 0 67436 0 -1 85952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_153_727
timestamp 1644511149
transform 1 0 67988 0 -1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_153_729
timestamp 1644511149
transform 1 0 68172 0 -1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_153_741
timestamp 1644511149
transform 1 0 69276 0 -1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_153_753
timestamp 1644511149
transform 1 0 70380 0 -1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_153_765
timestamp 1644511149
transform 1 0 71484 0 -1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_153_777
timestamp 1644511149
transform 1 0 72588 0 -1 85952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_153_783
timestamp 1644511149
transform 1 0 73140 0 -1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_153_785
timestamp 1644511149
transform 1 0 73324 0 -1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_153_797
timestamp 1644511149
transform 1 0 74428 0 -1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_153_809
timestamp 1644511149
transform 1 0 75532 0 -1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_153_821
timestamp 1644511149
transform 1 0 76636 0 -1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_153_833
timestamp 1644511149
transform 1 0 77740 0 -1 85952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_153_839
timestamp 1644511149
transform 1 0 78292 0 -1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_153_841
timestamp 1644511149
transform 1 0 78476 0 -1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_154_7
timestamp 1644511149
transform 1 0 1748 0 1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_154_19
timestamp 1644511149
transform 1 0 2852 0 1 85952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_154_27
timestamp 1644511149
transform 1 0 3588 0 1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_154_29
timestamp 1644511149
transform 1 0 3772 0 1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_154_41
timestamp 1644511149
transform 1 0 4876 0 1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_154_53
timestamp 1644511149
transform 1 0 5980 0 1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_154_65
timestamp 1644511149
transform 1 0 7084 0 1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_154_77
timestamp 1644511149
transform 1 0 8188 0 1 85952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_154_83
timestamp 1644511149
transform 1 0 8740 0 1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_154_85
timestamp 1644511149
transform 1 0 8924 0 1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_154_97
timestamp 1644511149
transform 1 0 10028 0 1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_154_109
timestamp 1644511149
transform 1 0 11132 0 1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_154_121
timestamp 1644511149
transform 1 0 12236 0 1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_154_133
timestamp 1644511149
transform 1 0 13340 0 1 85952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_154_139
timestamp 1644511149
transform 1 0 13892 0 1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_154_141
timestamp 1644511149
transform 1 0 14076 0 1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_154_153
timestamp 1644511149
transform 1 0 15180 0 1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_154_165
timestamp 1644511149
transform 1 0 16284 0 1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_154_177
timestamp 1644511149
transform 1 0 17388 0 1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_154_189
timestamp 1644511149
transform 1 0 18492 0 1 85952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_154_195
timestamp 1644511149
transform 1 0 19044 0 1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_154_197
timestamp 1644511149
transform 1 0 19228 0 1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_154_209
timestamp 1644511149
transform 1 0 20332 0 1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_154_221
timestamp 1644511149
transform 1 0 21436 0 1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_154_233
timestamp 1644511149
transform 1 0 22540 0 1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_154_245
timestamp 1644511149
transform 1 0 23644 0 1 85952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_154_251
timestamp 1644511149
transform 1 0 24196 0 1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_154_253
timestamp 1644511149
transform 1 0 24380 0 1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_154_265
timestamp 1644511149
transform 1 0 25484 0 1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_154_277
timestamp 1644511149
transform 1 0 26588 0 1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_154_289
timestamp 1644511149
transform 1 0 27692 0 1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_154_301
timestamp 1644511149
transform 1 0 28796 0 1 85952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_154_307
timestamp 1644511149
transform 1 0 29348 0 1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_154_309
timestamp 1644511149
transform 1 0 29532 0 1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_154_321
timestamp 1644511149
transform 1 0 30636 0 1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_154_333
timestamp 1644511149
transform 1 0 31740 0 1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_154_345
timestamp 1644511149
transform 1 0 32844 0 1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_154_357
timestamp 1644511149
transform 1 0 33948 0 1 85952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_154_363
timestamp 1644511149
transform 1 0 34500 0 1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_154_365
timestamp 1644511149
transform 1 0 34684 0 1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_154_377
timestamp 1644511149
transform 1 0 35788 0 1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_154_389
timestamp 1644511149
transform 1 0 36892 0 1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_154_401
timestamp 1644511149
transform 1 0 37996 0 1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_154_413
timestamp 1644511149
transform 1 0 39100 0 1 85952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_154_419
timestamp 1644511149
transform 1 0 39652 0 1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_154_421
timestamp 1644511149
transform 1 0 39836 0 1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_154_433
timestamp 1644511149
transform 1 0 40940 0 1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_154_445
timestamp 1644511149
transform 1 0 42044 0 1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_154_457
timestamp 1644511149
transform 1 0 43148 0 1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_154_469
timestamp 1644511149
transform 1 0 44252 0 1 85952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_154_475
timestamp 1644511149
transform 1 0 44804 0 1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_154_477
timestamp 1644511149
transform 1 0 44988 0 1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_154_489
timestamp 1644511149
transform 1 0 46092 0 1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_154_501
timestamp 1644511149
transform 1 0 47196 0 1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_154_513
timestamp 1644511149
transform 1 0 48300 0 1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_154_525
timestamp 1644511149
transform 1 0 49404 0 1 85952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_154_531
timestamp 1644511149
transform 1 0 49956 0 1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_154_533
timestamp 1644511149
transform 1 0 50140 0 1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_154_545
timestamp 1644511149
transform 1 0 51244 0 1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_154_557
timestamp 1644511149
transform 1 0 52348 0 1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_154_569
timestamp 1644511149
transform 1 0 53452 0 1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_154_581
timestamp 1644511149
transform 1 0 54556 0 1 85952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_154_587
timestamp 1644511149
transform 1 0 55108 0 1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_154_589
timestamp 1644511149
transform 1 0 55292 0 1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_154_601
timestamp 1644511149
transform 1 0 56396 0 1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_154_613
timestamp 1644511149
transform 1 0 57500 0 1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_154_625
timestamp 1644511149
transform 1 0 58604 0 1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_154_637
timestamp 1644511149
transform 1 0 59708 0 1 85952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_154_643
timestamp 1644511149
transform 1 0 60260 0 1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_154_645
timestamp 1644511149
transform 1 0 60444 0 1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_154_657
timestamp 1644511149
transform 1 0 61548 0 1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_154_669
timestamp 1644511149
transform 1 0 62652 0 1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_154_681
timestamp 1644511149
transform 1 0 63756 0 1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_154_693
timestamp 1644511149
transform 1 0 64860 0 1 85952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_154_699
timestamp 1644511149
transform 1 0 65412 0 1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_154_701
timestamp 1644511149
transform 1 0 65596 0 1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_154_713
timestamp 1644511149
transform 1 0 66700 0 1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_154_725
timestamp 1644511149
transform 1 0 67804 0 1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_154_737
timestamp 1644511149
transform 1 0 68908 0 1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_154_749
timestamp 1644511149
transform 1 0 70012 0 1 85952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_154_755
timestamp 1644511149
transform 1 0 70564 0 1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_154_757
timestamp 1644511149
transform 1 0 70748 0 1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_154_769
timestamp 1644511149
transform 1 0 71852 0 1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_154_781
timestamp 1644511149
transform 1 0 72956 0 1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_154_793
timestamp 1644511149
transform 1 0 74060 0 1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_154_805
timestamp 1644511149
transform 1 0 75164 0 1 85952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_154_811
timestamp 1644511149
transform 1 0 75716 0 1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_154_813
timestamp 1644511149
transform 1 0 75900 0 1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_154_825
timestamp 1644511149
transform 1 0 77004 0 1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_154_837
timestamp 1644511149
transform 1 0 78108 0 1 85952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_154_841
timestamp 1644511149
transform 1 0 78476 0 1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_155_3
timestamp 1644511149
transform 1 0 1380 0 -1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_155_15
timestamp 1644511149
transform 1 0 2484 0 -1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_155_27
timestamp 1644511149
transform 1 0 3588 0 -1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_155_39
timestamp 1644511149
transform 1 0 4692 0 -1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_155_51
timestamp 1644511149
transform 1 0 5796 0 -1 87040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_155_55
timestamp 1644511149
transform 1 0 6164 0 -1 87040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_155_57
timestamp 1644511149
transform 1 0 6348 0 -1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_155_69
timestamp 1644511149
transform 1 0 7452 0 -1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_155_81
timestamp 1644511149
transform 1 0 8556 0 -1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_155_93
timestamp 1644511149
transform 1 0 9660 0 -1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_155_105
timestamp 1644511149
transform 1 0 10764 0 -1 87040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_155_111
timestamp 1644511149
transform 1 0 11316 0 -1 87040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_155_113
timestamp 1644511149
transform 1 0 11500 0 -1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_155_125
timestamp 1644511149
transform 1 0 12604 0 -1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_155_137
timestamp 1644511149
transform 1 0 13708 0 -1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_155_149
timestamp 1644511149
transform 1 0 14812 0 -1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_155_161
timestamp 1644511149
transform 1 0 15916 0 -1 87040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_155_167
timestamp 1644511149
transform 1 0 16468 0 -1 87040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_155_169
timestamp 1644511149
transform 1 0 16652 0 -1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_155_181
timestamp 1644511149
transform 1 0 17756 0 -1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_155_193
timestamp 1644511149
transform 1 0 18860 0 -1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_155_205
timestamp 1644511149
transform 1 0 19964 0 -1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_155_217
timestamp 1644511149
transform 1 0 21068 0 -1 87040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_155_223
timestamp 1644511149
transform 1 0 21620 0 -1 87040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_155_225
timestamp 1644511149
transform 1 0 21804 0 -1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_155_237
timestamp 1644511149
transform 1 0 22908 0 -1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_155_249
timestamp 1644511149
transform 1 0 24012 0 -1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_155_261
timestamp 1644511149
transform 1 0 25116 0 -1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_155_273
timestamp 1644511149
transform 1 0 26220 0 -1 87040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_155_279
timestamp 1644511149
transform 1 0 26772 0 -1 87040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_155_281
timestamp 1644511149
transform 1 0 26956 0 -1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_155_293
timestamp 1644511149
transform 1 0 28060 0 -1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_155_305
timestamp 1644511149
transform 1 0 29164 0 -1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_155_317
timestamp 1644511149
transform 1 0 30268 0 -1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_155_329
timestamp 1644511149
transform 1 0 31372 0 -1 87040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_155_335
timestamp 1644511149
transform 1 0 31924 0 -1 87040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_155_337
timestamp 1644511149
transform 1 0 32108 0 -1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_155_349
timestamp 1644511149
transform 1 0 33212 0 -1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_155_361
timestamp 1644511149
transform 1 0 34316 0 -1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_155_373
timestamp 1644511149
transform 1 0 35420 0 -1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_155_385
timestamp 1644511149
transform 1 0 36524 0 -1 87040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_155_391
timestamp 1644511149
transform 1 0 37076 0 -1 87040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_155_393
timestamp 1644511149
transform 1 0 37260 0 -1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_155_405
timestamp 1644511149
transform 1 0 38364 0 -1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_155_417
timestamp 1644511149
transform 1 0 39468 0 -1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_155_429
timestamp 1644511149
transform 1 0 40572 0 -1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_155_441
timestamp 1644511149
transform 1 0 41676 0 -1 87040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_155_447
timestamp 1644511149
transform 1 0 42228 0 -1 87040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_155_449
timestamp 1644511149
transform 1 0 42412 0 -1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_155_461
timestamp 1644511149
transform 1 0 43516 0 -1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_155_473
timestamp 1644511149
transform 1 0 44620 0 -1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_155_485
timestamp 1644511149
transform 1 0 45724 0 -1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_155_497
timestamp 1644511149
transform 1 0 46828 0 -1 87040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_155_503
timestamp 1644511149
transform 1 0 47380 0 -1 87040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_155_505
timestamp 1644511149
transform 1 0 47564 0 -1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_155_517
timestamp 1644511149
transform 1 0 48668 0 -1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_155_529
timestamp 1644511149
transform 1 0 49772 0 -1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_155_541
timestamp 1644511149
transform 1 0 50876 0 -1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_155_553
timestamp 1644511149
transform 1 0 51980 0 -1 87040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_155_559
timestamp 1644511149
transform 1 0 52532 0 -1 87040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_155_561
timestamp 1644511149
transform 1 0 52716 0 -1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_155_573
timestamp 1644511149
transform 1 0 53820 0 -1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_155_585
timestamp 1644511149
transform 1 0 54924 0 -1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_155_597
timestamp 1644511149
transform 1 0 56028 0 -1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_155_609
timestamp 1644511149
transform 1 0 57132 0 -1 87040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_155_615
timestamp 1644511149
transform 1 0 57684 0 -1 87040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_155_617
timestamp 1644511149
transform 1 0 57868 0 -1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_155_629
timestamp 1644511149
transform 1 0 58972 0 -1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_155_641
timestamp 1644511149
transform 1 0 60076 0 -1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_155_653
timestamp 1644511149
transform 1 0 61180 0 -1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_155_665
timestamp 1644511149
transform 1 0 62284 0 -1 87040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_155_671
timestamp 1644511149
transform 1 0 62836 0 -1 87040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_155_673
timestamp 1644511149
transform 1 0 63020 0 -1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_155_685
timestamp 1644511149
transform 1 0 64124 0 -1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_155_697
timestamp 1644511149
transform 1 0 65228 0 -1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_155_709
timestamp 1644511149
transform 1 0 66332 0 -1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_155_721
timestamp 1644511149
transform 1 0 67436 0 -1 87040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_155_727
timestamp 1644511149
transform 1 0 67988 0 -1 87040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_155_729
timestamp 1644511149
transform 1 0 68172 0 -1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_155_741
timestamp 1644511149
transform 1 0 69276 0 -1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_155_753
timestamp 1644511149
transform 1 0 70380 0 -1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_155_765
timestamp 1644511149
transform 1 0 71484 0 -1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_155_777
timestamp 1644511149
transform 1 0 72588 0 -1 87040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_155_783
timestamp 1644511149
transform 1 0 73140 0 -1 87040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_155_785
timestamp 1644511149
transform 1 0 73324 0 -1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_155_797
timestamp 1644511149
transform 1 0 74428 0 -1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_155_809
timestamp 1644511149
transform 1 0 75532 0 -1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_155_821
timestamp 1644511149
transform 1 0 76636 0 -1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_155_833
timestamp 1644511149
transform 1 0 77740 0 -1 87040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_155_839
timestamp 1644511149
transform 1 0 78292 0 -1 87040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_155_841
timestamp 1644511149
transform 1 0 78476 0 -1 87040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_156_3
timestamp 1644511149
transform 1 0 1380 0 1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_156_15
timestamp 1644511149
transform 1 0 2484 0 1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_156_27
timestamp 1644511149
transform 1 0 3588 0 1 87040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_156_29
timestamp 1644511149
transform 1 0 3772 0 1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_156_41
timestamp 1644511149
transform 1 0 4876 0 1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_156_53
timestamp 1644511149
transform 1 0 5980 0 1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_156_65
timestamp 1644511149
transform 1 0 7084 0 1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_156_77
timestamp 1644511149
transform 1 0 8188 0 1 87040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_156_83
timestamp 1644511149
transform 1 0 8740 0 1 87040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_156_85
timestamp 1644511149
transform 1 0 8924 0 1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_156_97
timestamp 1644511149
transform 1 0 10028 0 1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_156_109
timestamp 1644511149
transform 1 0 11132 0 1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_156_121
timestamp 1644511149
transform 1 0 12236 0 1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_156_133
timestamp 1644511149
transform 1 0 13340 0 1 87040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_156_139
timestamp 1644511149
transform 1 0 13892 0 1 87040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_156_141
timestamp 1644511149
transform 1 0 14076 0 1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_156_153
timestamp 1644511149
transform 1 0 15180 0 1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_156_165
timestamp 1644511149
transform 1 0 16284 0 1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_156_177
timestamp 1644511149
transform 1 0 17388 0 1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_156_189
timestamp 1644511149
transform 1 0 18492 0 1 87040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_156_195
timestamp 1644511149
transform 1 0 19044 0 1 87040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_156_197
timestamp 1644511149
transform 1 0 19228 0 1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_156_209
timestamp 1644511149
transform 1 0 20332 0 1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_156_221
timestamp 1644511149
transform 1 0 21436 0 1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_156_233
timestamp 1644511149
transform 1 0 22540 0 1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_156_245
timestamp 1644511149
transform 1 0 23644 0 1 87040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_156_251
timestamp 1644511149
transform 1 0 24196 0 1 87040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_156_253
timestamp 1644511149
transform 1 0 24380 0 1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_156_265
timestamp 1644511149
transform 1 0 25484 0 1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_156_277
timestamp 1644511149
transform 1 0 26588 0 1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_156_289
timestamp 1644511149
transform 1 0 27692 0 1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_156_301
timestamp 1644511149
transform 1 0 28796 0 1 87040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_156_307
timestamp 1644511149
transform 1 0 29348 0 1 87040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_156_309
timestamp 1644511149
transform 1 0 29532 0 1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_156_321
timestamp 1644511149
transform 1 0 30636 0 1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_156_333
timestamp 1644511149
transform 1 0 31740 0 1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_156_345
timestamp 1644511149
transform 1 0 32844 0 1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_156_357
timestamp 1644511149
transform 1 0 33948 0 1 87040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_156_363
timestamp 1644511149
transform 1 0 34500 0 1 87040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_156_365
timestamp 1644511149
transform 1 0 34684 0 1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_156_377
timestamp 1644511149
transform 1 0 35788 0 1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_156_389
timestamp 1644511149
transform 1 0 36892 0 1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_156_401
timestamp 1644511149
transform 1 0 37996 0 1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_156_413
timestamp 1644511149
transform 1 0 39100 0 1 87040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_156_419
timestamp 1644511149
transform 1 0 39652 0 1 87040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_156_421
timestamp 1644511149
transform 1 0 39836 0 1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_156_433
timestamp 1644511149
transform 1 0 40940 0 1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_156_445
timestamp 1644511149
transform 1 0 42044 0 1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_156_457
timestamp 1644511149
transform 1 0 43148 0 1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_156_469
timestamp 1644511149
transform 1 0 44252 0 1 87040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_156_475
timestamp 1644511149
transform 1 0 44804 0 1 87040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_156_477
timestamp 1644511149
transform 1 0 44988 0 1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_156_489
timestamp 1644511149
transform 1 0 46092 0 1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_156_501
timestamp 1644511149
transform 1 0 47196 0 1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_156_513
timestamp 1644511149
transform 1 0 48300 0 1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_156_525
timestamp 1644511149
transform 1 0 49404 0 1 87040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_156_531
timestamp 1644511149
transform 1 0 49956 0 1 87040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_156_533
timestamp 1644511149
transform 1 0 50140 0 1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_156_545
timestamp 1644511149
transform 1 0 51244 0 1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_156_557
timestamp 1644511149
transform 1 0 52348 0 1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_156_569
timestamp 1644511149
transform 1 0 53452 0 1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_156_581
timestamp 1644511149
transform 1 0 54556 0 1 87040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_156_587
timestamp 1644511149
transform 1 0 55108 0 1 87040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_156_589
timestamp 1644511149
transform 1 0 55292 0 1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_156_601
timestamp 1644511149
transform 1 0 56396 0 1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_156_613
timestamp 1644511149
transform 1 0 57500 0 1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_156_625
timestamp 1644511149
transform 1 0 58604 0 1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_156_637
timestamp 1644511149
transform 1 0 59708 0 1 87040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_156_643
timestamp 1644511149
transform 1 0 60260 0 1 87040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_156_645
timestamp 1644511149
transform 1 0 60444 0 1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_156_657
timestamp 1644511149
transform 1 0 61548 0 1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_156_669
timestamp 1644511149
transform 1 0 62652 0 1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_156_681
timestamp 1644511149
transform 1 0 63756 0 1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_156_693
timestamp 1644511149
transform 1 0 64860 0 1 87040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_156_699
timestamp 1644511149
transform 1 0 65412 0 1 87040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_156_701
timestamp 1644511149
transform 1 0 65596 0 1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_156_713
timestamp 1644511149
transform 1 0 66700 0 1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_156_725
timestamp 1644511149
transform 1 0 67804 0 1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_156_737
timestamp 1644511149
transform 1 0 68908 0 1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_156_749
timestamp 1644511149
transform 1 0 70012 0 1 87040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_156_755
timestamp 1644511149
transform 1 0 70564 0 1 87040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_156_757
timestamp 1644511149
transform 1 0 70748 0 1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_156_769
timestamp 1644511149
transform 1 0 71852 0 1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_156_781
timestamp 1644511149
transform 1 0 72956 0 1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_156_793
timestamp 1644511149
transform 1 0 74060 0 1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_156_805
timestamp 1644511149
transform 1 0 75164 0 1 87040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_156_811
timestamp 1644511149
transform 1 0 75716 0 1 87040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_156_813
timestamp 1644511149
transform 1 0 75900 0 1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_156_825
timestamp 1644511149
transform 1 0 77004 0 1 87040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_156_831
timestamp 1644511149
transform 1 0 77556 0 1 87040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_156_838
timestamp 1644511149
transform 1 0 78200 0 1 87040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_157_3
timestamp 1644511149
transform 1 0 1380 0 -1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_157_15
timestamp 1644511149
transform 1 0 2484 0 -1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_157_27
timestamp 1644511149
transform 1 0 3588 0 -1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_157_39
timestamp 1644511149
transform 1 0 4692 0 -1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_157_51
timestamp 1644511149
transform 1 0 5796 0 -1 88128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_157_55
timestamp 1644511149
transform 1 0 6164 0 -1 88128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_157_57
timestamp 1644511149
transform 1 0 6348 0 -1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_157_69
timestamp 1644511149
transform 1 0 7452 0 -1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_157_81
timestamp 1644511149
transform 1 0 8556 0 -1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_157_93
timestamp 1644511149
transform 1 0 9660 0 -1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_157_105
timestamp 1644511149
transform 1 0 10764 0 -1 88128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_157_111
timestamp 1644511149
transform 1 0 11316 0 -1 88128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_157_113
timestamp 1644511149
transform 1 0 11500 0 -1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_157_125
timestamp 1644511149
transform 1 0 12604 0 -1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_157_137
timestamp 1644511149
transform 1 0 13708 0 -1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_157_149
timestamp 1644511149
transform 1 0 14812 0 -1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_157_161
timestamp 1644511149
transform 1 0 15916 0 -1 88128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_157_167
timestamp 1644511149
transform 1 0 16468 0 -1 88128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_157_169
timestamp 1644511149
transform 1 0 16652 0 -1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_157_181
timestamp 1644511149
transform 1 0 17756 0 -1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_157_193
timestamp 1644511149
transform 1 0 18860 0 -1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_157_205
timestamp 1644511149
transform 1 0 19964 0 -1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_157_217
timestamp 1644511149
transform 1 0 21068 0 -1 88128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_157_223
timestamp 1644511149
transform 1 0 21620 0 -1 88128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_157_225
timestamp 1644511149
transform 1 0 21804 0 -1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_157_237
timestamp 1644511149
transform 1 0 22908 0 -1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_157_249
timestamp 1644511149
transform 1 0 24012 0 -1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_157_261
timestamp 1644511149
transform 1 0 25116 0 -1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_157_273
timestamp 1644511149
transform 1 0 26220 0 -1 88128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_157_279
timestamp 1644511149
transform 1 0 26772 0 -1 88128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_157_281
timestamp 1644511149
transform 1 0 26956 0 -1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_157_293
timestamp 1644511149
transform 1 0 28060 0 -1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_157_305
timestamp 1644511149
transform 1 0 29164 0 -1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_157_317
timestamp 1644511149
transform 1 0 30268 0 -1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_157_329
timestamp 1644511149
transform 1 0 31372 0 -1 88128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_157_335
timestamp 1644511149
transform 1 0 31924 0 -1 88128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_157_337
timestamp 1644511149
transform 1 0 32108 0 -1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_157_349
timestamp 1644511149
transform 1 0 33212 0 -1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_157_361
timestamp 1644511149
transform 1 0 34316 0 -1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_157_373
timestamp 1644511149
transform 1 0 35420 0 -1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_157_385
timestamp 1644511149
transform 1 0 36524 0 -1 88128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_157_391
timestamp 1644511149
transform 1 0 37076 0 -1 88128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_157_393
timestamp 1644511149
transform 1 0 37260 0 -1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_157_405
timestamp 1644511149
transform 1 0 38364 0 -1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_157_417
timestamp 1644511149
transform 1 0 39468 0 -1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_157_429
timestamp 1644511149
transform 1 0 40572 0 -1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_157_441
timestamp 1644511149
transform 1 0 41676 0 -1 88128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_157_447
timestamp 1644511149
transform 1 0 42228 0 -1 88128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_157_449
timestamp 1644511149
transform 1 0 42412 0 -1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_157_461
timestamp 1644511149
transform 1 0 43516 0 -1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_157_473
timestamp 1644511149
transform 1 0 44620 0 -1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_157_485
timestamp 1644511149
transform 1 0 45724 0 -1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_157_497
timestamp 1644511149
transform 1 0 46828 0 -1 88128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_157_503
timestamp 1644511149
transform 1 0 47380 0 -1 88128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_157_505
timestamp 1644511149
transform 1 0 47564 0 -1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_157_517
timestamp 1644511149
transform 1 0 48668 0 -1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_157_529
timestamp 1644511149
transform 1 0 49772 0 -1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_157_541
timestamp 1644511149
transform 1 0 50876 0 -1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_157_553
timestamp 1644511149
transform 1 0 51980 0 -1 88128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_157_559
timestamp 1644511149
transform 1 0 52532 0 -1 88128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_157_561
timestamp 1644511149
transform 1 0 52716 0 -1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_157_573
timestamp 1644511149
transform 1 0 53820 0 -1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_157_585
timestamp 1644511149
transform 1 0 54924 0 -1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_157_597
timestamp 1644511149
transform 1 0 56028 0 -1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_157_609
timestamp 1644511149
transform 1 0 57132 0 -1 88128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_157_615
timestamp 1644511149
transform 1 0 57684 0 -1 88128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_157_617
timestamp 1644511149
transform 1 0 57868 0 -1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_157_629
timestamp 1644511149
transform 1 0 58972 0 -1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_157_641
timestamp 1644511149
transform 1 0 60076 0 -1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_157_653
timestamp 1644511149
transform 1 0 61180 0 -1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_157_665
timestamp 1644511149
transform 1 0 62284 0 -1 88128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_157_671
timestamp 1644511149
transform 1 0 62836 0 -1 88128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_157_673
timestamp 1644511149
transform 1 0 63020 0 -1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_157_685
timestamp 1644511149
transform 1 0 64124 0 -1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_157_697
timestamp 1644511149
transform 1 0 65228 0 -1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_157_709
timestamp 1644511149
transform 1 0 66332 0 -1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_157_721
timestamp 1644511149
transform 1 0 67436 0 -1 88128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_157_727
timestamp 1644511149
transform 1 0 67988 0 -1 88128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_157_729
timestamp 1644511149
transform 1 0 68172 0 -1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_157_741
timestamp 1644511149
transform 1 0 69276 0 -1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_157_753
timestamp 1644511149
transform 1 0 70380 0 -1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_157_765
timestamp 1644511149
transform 1 0 71484 0 -1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_157_777
timestamp 1644511149
transform 1 0 72588 0 -1 88128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_157_783
timestamp 1644511149
transform 1 0 73140 0 -1 88128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_157_785
timestamp 1644511149
transform 1 0 73324 0 -1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_157_797
timestamp 1644511149
transform 1 0 74428 0 -1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_157_809
timestamp 1644511149
transform 1 0 75532 0 -1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_157_821
timestamp 1644511149
transform 1 0 76636 0 -1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_157_833
timestamp 1644511149
transform 1 0 77740 0 -1 88128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_157_839
timestamp 1644511149
transform 1 0 78292 0 -1 88128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_157_841
timestamp 1644511149
transform 1 0 78476 0 -1 88128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_158_3
timestamp 1644511149
transform 1 0 1380 0 1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_158_15
timestamp 1644511149
transform 1 0 2484 0 1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_158_27
timestamp 1644511149
transform 1 0 3588 0 1 88128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_158_29
timestamp 1644511149
transform 1 0 3772 0 1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_158_41
timestamp 1644511149
transform 1 0 4876 0 1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_158_53
timestamp 1644511149
transform 1 0 5980 0 1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_158_65
timestamp 1644511149
transform 1 0 7084 0 1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_158_77
timestamp 1644511149
transform 1 0 8188 0 1 88128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_158_83
timestamp 1644511149
transform 1 0 8740 0 1 88128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_158_85
timestamp 1644511149
transform 1 0 8924 0 1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_158_97
timestamp 1644511149
transform 1 0 10028 0 1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_158_109
timestamp 1644511149
transform 1 0 11132 0 1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_158_121
timestamp 1644511149
transform 1 0 12236 0 1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_158_133
timestamp 1644511149
transform 1 0 13340 0 1 88128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_158_139
timestamp 1644511149
transform 1 0 13892 0 1 88128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_158_141
timestamp 1644511149
transform 1 0 14076 0 1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_158_153
timestamp 1644511149
transform 1 0 15180 0 1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_158_165
timestamp 1644511149
transform 1 0 16284 0 1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_158_177
timestamp 1644511149
transform 1 0 17388 0 1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_158_189
timestamp 1644511149
transform 1 0 18492 0 1 88128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_158_195
timestamp 1644511149
transform 1 0 19044 0 1 88128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_158_197
timestamp 1644511149
transform 1 0 19228 0 1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_158_209
timestamp 1644511149
transform 1 0 20332 0 1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_158_221
timestamp 1644511149
transform 1 0 21436 0 1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_158_233
timestamp 1644511149
transform 1 0 22540 0 1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_158_245
timestamp 1644511149
transform 1 0 23644 0 1 88128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_158_251
timestamp 1644511149
transform 1 0 24196 0 1 88128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_158_253
timestamp 1644511149
transform 1 0 24380 0 1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_158_265
timestamp 1644511149
transform 1 0 25484 0 1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_158_277
timestamp 1644511149
transform 1 0 26588 0 1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_158_289
timestamp 1644511149
transform 1 0 27692 0 1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_158_301
timestamp 1644511149
transform 1 0 28796 0 1 88128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_158_307
timestamp 1644511149
transform 1 0 29348 0 1 88128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_158_309
timestamp 1644511149
transform 1 0 29532 0 1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_158_321
timestamp 1644511149
transform 1 0 30636 0 1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_158_333
timestamp 1644511149
transform 1 0 31740 0 1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_158_345
timestamp 1644511149
transform 1 0 32844 0 1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_158_357
timestamp 1644511149
transform 1 0 33948 0 1 88128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_158_363
timestamp 1644511149
transform 1 0 34500 0 1 88128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_158_365
timestamp 1644511149
transform 1 0 34684 0 1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_158_377
timestamp 1644511149
transform 1 0 35788 0 1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_158_389
timestamp 1644511149
transform 1 0 36892 0 1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_158_401
timestamp 1644511149
transform 1 0 37996 0 1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_158_413
timestamp 1644511149
transform 1 0 39100 0 1 88128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_158_419
timestamp 1644511149
transform 1 0 39652 0 1 88128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_158_421
timestamp 1644511149
transform 1 0 39836 0 1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_158_433
timestamp 1644511149
transform 1 0 40940 0 1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_158_445
timestamp 1644511149
transform 1 0 42044 0 1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_158_457
timestamp 1644511149
transform 1 0 43148 0 1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_158_469
timestamp 1644511149
transform 1 0 44252 0 1 88128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_158_475
timestamp 1644511149
transform 1 0 44804 0 1 88128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_158_477
timestamp 1644511149
transform 1 0 44988 0 1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_158_489
timestamp 1644511149
transform 1 0 46092 0 1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_158_501
timestamp 1644511149
transform 1 0 47196 0 1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_158_513
timestamp 1644511149
transform 1 0 48300 0 1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_158_525
timestamp 1644511149
transform 1 0 49404 0 1 88128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_158_531
timestamp 1644511149
transform 1 0 49956 0 1 88128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_158_533
timestamp 1644511149
transform 1 0 50140 0 1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_158_545
timestamp 1644511149
transform 1 0 51244 0 1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_158_557
timestamp 1644511149
transform 1 0 52348 0 1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_158_569
timestamp 1644511149
transform 1 0 53452 0 1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_158_581
timestamp 1644511149
transform 1 0 54556 0 1 88128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_158_587
timestamp 1644511149
transform 1 0 55108 0 1 88128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_158_589
timestamp 1644511149
transform 1 0 55292 0 1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_158_601
timestamp 1644511149
transform 1 0 56396 0 1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_158_613
timestamp 1644511149
transform 1 0 57500 0 1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_158_625
timestamp 1644511149
transform 1 0 58604 0 1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_158_637
timestamp 1644511149
transform 1 0 59708 0 1 88128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_158_643
timestamp 1644511149
transform 1 0 60260 0 1 88128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_158_645
timestamp 1644511149
transform 1 0 60444 0 1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_158_657
timestamp 1644511149
transform 1 0 61548 0 1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_158_669
timestamp 1644511149
transform 1 0 62652 0 1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_158_681
timestamp 1644511149
transform 1 0 63756 0 1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_158_693
timestamp 1644511149
transform 1 0 64860 0 1 88128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_158_699
timestamp 1644511149
transform 1 0 65412 0 1 88128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_158_701
timestamp 1644511149
transform 1 0 65596 0 1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_158_713
timestamp 1644511149
transform 1 0 66700 0 1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_158_725
timestamp 1644511149
transform 1 0 67804 0 1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_158_737
timestamp 1644511149
transform 1 0 68908 0 1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_158_749
timestamp 1644511149
transform 1 0 70012 0 1 88128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_158_755
timestamp 1644511149
transform 1 0 70564 0 1 88128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_158_757
timestamp 1644511149
transform 1 0 70748 0 1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_158_769
timestamp 1644511149
transform 1 0 71852 0 1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_158_781
timestamp 1644511149
transform 1 0 72956 0 1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_158_793
timestamp 1644511149
transform 1 0 74060 0 1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_158_805
timestamp 1644511149
transform 1 0 75164 0 1 88128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_158_811
timestamp 1644511149
transform 1 0 75716 0 1 88128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_158_813
timestamp 1644511149
transform 1 0 75900 0 1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_158_825
timestamp 1644511149
transform 1 0 77004 0 1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_158_837
timestamp 1644511149
transform 1 0 78108 0 1 88128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_158_841
timestamp 1644511149
transform 1 0 78476 0 1 88128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_159_3
timestamp 1644511149
transform 1 0 1380 0 -1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_159_15
timestamp 1644511149
transform 1 0 2484 0 -1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_159_27
timestamp 1644511149
transform 1 0 3588 0 -1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_159_39
timestamp 1644511149
transform 1 0 4692 0 -1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_159_51
timestamp 1644511149
transform 1 0 5796 0 -1 89216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_159_55
timestamp 1644511149
transform 1 0 6164 0 -1 89216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_159_57
timestamp 1644511149
transform 1 0 6348 0 -1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_159_69
timestamp 1644511149
transform 1 0 7452 0 -1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_159_81
timestamp 1644511149
transform 1 0 8556 0 -1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_159_93
timestamp 1644511149
transform 1 0 9660 0 -1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_159_105
timestamp 1644511149
transform 1 0 10764 0 -1 89216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_159_111
timestamp 1644511149
transform 1 0 11316 0 -1 89216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_159_113
timestamp 1644511149
transform 1 0 11500 0 -1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_159_125
timestamp 1644511149
transform 1 0 12604 0 -1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_159_137
timestamp 1644511149
transform 1 0 13708 0 -1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_159_149
timestamp 1644511149
transform 1 0 14812 0 -1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_159_161
timestamp 1644511149
transform 1 0 15916 0 -1 89216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_159_167
timestamp 1644511149
transform 1 0 16468 0 -1 89216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_159_169
timestamp 1644511149
transform 1 0 16652 0 -1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_159_181
timestamp 1644511149
transform 1 0 17756 0 -1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_159_193
timestamp 1644511149
transform 1 0 18860 0 -1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_159_205
timestamp 1644511149
transform 1 0 19964 0 -1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_159_217
timestamp 1644511149
transform 1 0 21068 0 -1 89216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_159_223
timestamp 1644511149
transform 1 0 21620 0 -1 89216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_159_225
timestamp 1644511149
transform 1 0 21804 0 -1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_159_237
timestamp 1644511149
transform 1 0 22908 0 -1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_159_249
timestamp 1644511149
transform 1 0 24012 0 -1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_159_261
timestamp 1644511149
transform 1 0 25116 0 -1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_159_273
timestamp 1644511149
transform 1 0 26220 0 -1 89216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_159_279
timestamp 1644511149
transform 1 0 26772 0 -1 89216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_159_281
timestamp 1644511149
transform 1 0 26956 0 -1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_159_293
timestamp 1644511149
transform 1 0 28060 0 -1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_159_305
timestamp 1644511149
transform 1 0 29164 0 -1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_159_317
timestamp 1644511149
transform 1 0 30268 0 -1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_159_329
timestamp 1644511149
transform 1 0 31372 0 -1 89216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_159_335
timestamp 1644511149
transform 1 0 31924 0 -1 89216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_159_337
timestamp 1644511149
transform 1 0 32108 0 -1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_159_349
timestamp 1644511149
transform 1 0 33212 0 -1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_159_361
timestamp 1644511149
transform 1 0 34316 0 -1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_159_373
timestamp 1644511149
transform 1 0 35420 0 -1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_159_385
timestamp 1644511149
transform 1 0 36524 0 -1 89216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_159_391
timestamp 1644511149
transform 1 0 37076 0 -1 89216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_159_393
timestamp 1644511149
transform 1 0 37260 0 -1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_159_405
timestamp 1644511149
transform 1 0 38364 0 -1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_159_417
timestamp 1644511149
transform 1 0 39468 0 -1 89216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_159_427
timestamp 1644511149
transform 1 0 40388 0 -1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_159_439
timestamp 1644511149
transform 1 0 41492 0 -1 89216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_159_447
timestamp 1644511149
transform 1 0 42228 0 -1 89216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_159_449
timestamp 1644511149
transform 1 0 42412 0 -1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_159_461
timestamp 1644511149
transform 1 0 43516 0 -1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_159_473
timestamp 1644511149
transform 1 0 44620 0 -1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_159_485
timestamp 1644511149
transform 1 0 45724 0 -1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_159_497
timestamp 1644511149
transform 1 0 46828 0 -1 89216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_159_503
timestamp 1644511149
transform 1 0 47380 0 -1 89216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_159_505
timestamp 1644511149
transform 1 0 47564 0 -1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_159_517
timestamp 1644511149
transform 1 0 48668 0 -1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_159_529
timestamp 1644511149
transform 1 0 49772 0 -1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_159_541
timestamp 1644511149
transform 1 0 50876 0 -1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_159_553
timestamp 1644511149
transform 1 0 51980 0 -1 89216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_159_559
timestamp 1644511149
transform 1 0 52532 0 -1 89216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_159_561
timestamp 1644511149
transform 1 0 52716 0 -1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_159_573
timestamp 1644511149
transform 1 0 53820 0 -1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_159_585
timestamp 1644511149
transform 1 0 54924 0 -1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_159_597
timestamp 1644511149
transform 1 0 56028 0 -1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_159_609
timestamp 1644511149
transform 1 0 57132 0 -1 89216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_159_615
timestamp 1644511149
transform 1 0 57684 0 -1 89216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_159_617
timestamp 1644511149
transform 1 0 57868 0 -1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_159_629
timestamp 1644511149
transform 1 0 58972 0 -1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_159_641
timestamp 1644511149
transform 1 0 60076 0 -1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_159_653
timestamp 1644511149
transform 1 0 61180 0 -1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_159_665
timestamp 1644511149
transform 1 0 62284 0 -1 89216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_159_671
timestamp 1644511149
transform 1 0 62836 0 -1 89216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_159_673
timestamp 1644511149
transform 1 0 63020 0 -1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_159_685
timestamp 1644511149
transform 1 0 64124 0 -1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_159_697
timestamp 1644511149
transform 1 0 65228 0 -1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_159_709
timestamp 1644511149
transform 1 0 66332 0 -1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_159_721
timestamp 1644511149
transform 1 0 67436 0 -1 89216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_159_727
timestamp 1644511149
transform 1 0 67988 0 -1 89216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_159_729
timestamp 1644511149
transform 1 0 68172 0 -1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_159_741
timestamp 1644511149
transform 1 0 69276 0 -1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_159_753
timestamp 1644511149
transform 1 0 70380 0 -1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_159_765
timestamp 1644511149
transform 1 0 71484 0 -1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_159_777
timestamp 1644511149
transform 1 0 72588 0 -1 89216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_159_783
timestamp 1644511149
transform 1 0 73140 0 -1 89216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_159_785
timestamp 1644511149
transform 1 0 73324 0 -1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_159_797
timestamp 1644511149
transform 1 0 74428 0 -1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_159_809
timestamp 1644511149
transform 1 0 75532 0 -1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_159_821
timestamp 1644511149
transform 1 0 76636 0 -1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_159_833
timestamp 1644511149
transform 1 0 77740 0 -1 89216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_159_839
timestamp 1644511149
transform 1 0 78292 0 -1 89216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_159_841
timestamp 1644511149
transform 1 0 78476 0 -1 89216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_160_3
timestamp 1644511149
transform 1 0 1380 0 1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_160_15
timestamp 1644511149
transform 1 0 2484 0 1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_160_27
timestamp 1644511149
transform 1 0 3588 0 1 89216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_160_29
timestamp 1644511149
transform 1 0 3772 0 1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_160_41
timestamp 1644511149
transform 1 0 4876 0 1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_160_53
timestamp 1644511149
transform 1 0 5980 0 1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_160_65
timestamp 1644511149
transform 1 0 7084 0 1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_160_77
timestamp 1644511149
transform 1 0 8188 0 1 89216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_160_83
timestamp 1644511149
transform 1 0 8740 0 1 89216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_160_85
timestamp 1644511149
transform 1 0 8924 0 1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_160_97
timestamp 1644511149
transform 1 0 10028 0 1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_160_109
timestamp 1644511149
transform 1 0 11132 0 1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_160_121
timestamp 1644511149
transform 1 0 12236 0 1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_160_133
timestamp 1644511149
transform 1 0 13340 0 1 89216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_160_139
timestamp 1644511149
transform 1 0 13892 0 1 89216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_160_141
timestamp 1644511149
transform 1 0 14076 0 1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_160_153
timestamp 1644511149
transform 1 0 15180 0 1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_160_165
timestamp 1644511149
transform 1 0 16284 0 1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_160_177
timestamp 1644511149
transform 1 0 17388 0 1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_160_189
timestamp 1644511149
transform 1 0 18492 0 1 89216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_160_195
timestamp 1644511149
transform 1 0 19044 0 1 89216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_160_197
timestamp 1644511149
transform 1 0 19228 0 1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_160_209
timestamp 1644511149
transform 1 0 20332 0 1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_160_221
timestamp 1644511149
transform 1 0 21436 0 1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_160_233
timestamp 1644511149
transform 1 0 22540 0 1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_160_245
timestamp 1644511149
transform 1 0 23644 0 1 89216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_160_251
timestamp 1644511149
transform 1 0 24196 0 1 89216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_160_253
timestamp 1644511149
transform 1 0 24380 0 1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_160_265
timestamp 1644511149
transform 1 0 25484 0 1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_160_277
timestamp 1644511149
transform 1 0 26588 0 1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_160_289
timestamp 1644511149
transform 1 0 27692 0 1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_160_301
timestamp 1644511149
transform 1 0 28796 0 1 89216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_160_307
timestamp 1644511149
transform 1 0 29348 0 1 89216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_160_309
timestamp 1644511149
transform 1 0 29532 0 1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_160_321
timestamp 1644511149
transform 1 0 30636 0 1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_160_333
timestamp 1644511149
transform 1 0 31740 0 1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_160_345
timestamp 1644511149
transform 1 0 32844 0 1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_160_357
timestamp 1644511149
transform 1 0 33948 0 1 89216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_160_363
timestamp 1644511149
transform 1 0 34500 0 1 89216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_160_365
timestamp 1644511149
transform 1 0 34684 0 1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_160_377
timestamp 1644511149
transform 1 0 35788 0 1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_160_389
timestamp 1644511149
transform 1 0 36892 0 1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_160_401
timestamp 1644511149
transform 1 0 37996 0 1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_160_413
timestamp 1644511149
transform 1 0 39100 0 1 89216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_160_419
timestamp 1644511149
transform 1 0 39652 0 1 89216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_160_421
timestamp 1644511149
transform 1 0 39836 0 1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_160_433
timestamp 1644511149
transform 1 0 40940 0 1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_160_445
timestamp 1644511149
transform 1 0 42044 0 1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_160_457
timestamp 1644511149
transform 1 0 43148 0 1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_160_469
timestamp 1644511149
transform 1 0 44252 0 1 89216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_160_475
timestamp 1644511149
transform 1 0 44804 0 1 89216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_160_477
timestamp 1644511149
transform 1 0 44988 0 1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_160_489
timestamp 1644511149
transform 1 0 46092 0 1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_160_501
timestamp 1644511149
transform 1 0 47196 0 1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_160_513
timestamp 1644511149
transform 1 0 48300 0 1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_160_525
timestamp 1644511149
transform 1 0 49404 0 1 89216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_160_531
timestamp 1644511149
transform 1 0 49956 0 1 89216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_160_533
timestamp 1644511149
transform 1 0 50140 0 1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_160_545
timestamp 1644511149
transform 1 0 51244 0 1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_160_557
timestamp 1644511149
transform 1 0 52348 0 1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_160_569
timestamp 1644511149
transform 1 0 53452 0 1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_160_581
timestamp 1644511149
transform 1 0 54556 0 1 89216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_160_587
timestamp 1644511149
transform 1 0 55108 0 1 89216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_160_589
timestamp 1644511149
transform 1 0 55292 0 1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_160_601
timestamp 1644511149
transform 1 0 56396 0 1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_160_613
timestamp 1644511149
transform 1 0 57500 0 1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_160_625
timestamp 1644511149
transform 1 0 58604 0 1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_160_637
timestamp 1644511149
transform 1 0 59708 0 1 89216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_160_643
timestamp 1644511149
transform 1 0 60260 0 1 89216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_160_645
timestamp 1644511149
transform 1 0 60444 0 1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_160_657
timestamp 1644511149
transform 1 0 61548 0 1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_160_669
timestamp 1644511149
transform 1 0 62652 0 1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_160_681
timestamp 1644511149
transform 1 0 63756 0 1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_160_693
timestamp 1644511149
transform 1 0 64860 0 1 89216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_160_699
timestamp 1644511149
transform 1 0 65412 0 1 89216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_160_701
timestamp 1644511149
transform 1 0 65596 0 1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_160_713
timestamp 1644511149
transform 1 0 66700 0 1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_160_725
timestamp 1644511149
transform 1 0 67804 0 1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_160_737
timestamp 1644511149
transform 1 0 68908 0 1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_160_749
timestamp 1644511149
transform 1 0 70012 0 1 89216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_160_755
timestamp 1644511149
transform 1 0 70564 0 1 89216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_160_757
timestamp 1644511149
transform 1 0 70748 0 1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_160_769
timestamp 1644511149
transform 1 0 71852 0 1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_160_781
timestamp 1644511149
transform 1 0 72956 0 1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_160_793
timestamp 1644511149
transform 1 0 74060 0 1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_160_805
timestamp 1644511149
transform 1 0 75164 0 1 89216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_160_811
timestamp 1644511149
transform 1 0 75716 0 1 89216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_160_813
timestamp 1644511149
transform 1 0 75900 0 1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_160_825
timestamp 1644511149
transform 1 0 77004 0 1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_160_837
timestamp 1644511149
transform 1 0 78108 0 1 89216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_160_841
timestamp 1644511149
transform 1 0 78476 0 1 89216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_161_12
timestamp 1644511149
transform 1 0 2208 0 -1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_161_24
timestamp 1644511149
transform 1 0 3312 0 -1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_161_36
timestamp 1644511149
transform 1 0 4416 0 -1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_161_48
timestamp 1644511149
transform 1 0 5520 0 -1 90304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_161_57
timestamp 1644511149
transform 1 0 6348 0 -1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_161_69
timestamp 1644511149
transform 1 0 7452 0 -1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_161_81
timestamp 1644511149
transform 1 0 8556 0 -1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_161_93
timestamp 1644511149
transform 1 0 9660 0 -1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_161_105
timestamp 1644511149
transform 1 0 10764 0 -1 90304
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_161_111
timestamp 1644511149
transform 1 0 11316 0 -1 90304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_161_113
timestamp 1644511149
transform 1 0 11500 0 -1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_161_125
timestamp 1644511149
transform 1 0 12604 0 -1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_161_137
timestamp 1644511149
transform 1 0 13708 0 -1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_161_149
timestamp 1644511149
transform 1 0 14812 0 -1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_161_161
timestamp 1644511149
transform 1 0 15916 0 -1 90304
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_161_167
timestamp 1644511149
transform 1 0 16468 0 -1 90304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_161_169
timestamp 1644511149
transform 1 0 16652 0 -1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_161_181
timestamp 1644511149
transform 1 0 17756 0 -1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_161_193
timestamp 1644511149
transform 1 0 18860 0 -1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_161_205
timestamp 1644511149
transform 1 0 19964 0 -1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_161_217
timestamp 1644511149
transform 1 0 21068 0 -1 90304
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_161_223
timestamp 1644511149
transform 1 0 21620 0 -1 90304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_161_225
timestamp 1644511149
transform 1 0 21804 0 -1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_161_237
timestamp 1644511149
transform 1 0 22908 0 -1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_161_249
timestamp 1644511149
transform 1 0 24012 0 -1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_161_261
timestamp 1644511149
transform 1 0 25116 0 -1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_161_273
timestamp 1644511149
transform 1 0 26220 0 -1 90304
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_161_279
timestamp 1644511149
transform 1 0 26772 0 -1 90304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_161_281
timestamp 1644511149
transform 1 0 26956 0 -1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_161_293
timestamp 1644511149
transform 1 0 28060 0 -1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_161_305
timestamp 1644511149
transform 1 0 29164 0 -1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_161_317
timestamp 1644511149
transform 1 0 30268 0 -1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_161_329
timestamp 1644511149
transform 1 0 31372 0 -1 90304
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_161_335
timestamp 1644511149
transform 1 0 31924 0 -1 90304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_161_337
timestamp 1644511149
transform 1 0 32108 0 -1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_161_349
timestamp 1644511149
transform 1 0 33212 0 -1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_161_361
timestamp 1644511149
transform 1 0 34316 0 -1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_161_373
timestamp 1644511149
transform 1 0 35420 0 -1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_161_385
timestamp 1644511149
transform 1 0 36524 0 -1 90304
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_161_391
timestamp 1644511149
transform 1 0 37076 0 -1 90304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_161_393
timestamp 1644511149
transform 1 0 37260 0 -1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_161_405
timestamp 1644511149
transform 1 0 38364 0 -1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_161_417
timestamp 1644511149
transform 1 0 39468 0 -1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_161_429
timestamp 1644511149
transform 1 0 40572 0 -1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_161_441
timestamp 1644511149
transform 1 0 41676 0 -1 90304
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_161_447
timestamp 1644511149
transform 1 0 42228 0 -1 90304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_161_449
timestamp 1644511149
transform 1 0 42412 0 -1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_161_461
timestamp 1644511149
transform 1 0 43516 0 -1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_161_473
timestamp 1644511149
transform 1 0 44620 0 -1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_161_485
timestamp 1644511149
transform 1 0 45724 0 -1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_161_497
timestamp 1644511149
transform 1 0 46828 0 -1 90304
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_161_503
timestamp 1644511149
transform 1 0 47380 0 -1 90304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_161_505
timestamp 1644511149
transform 1 0 47564 0 -1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_161_517
timestamp 1644511149
transform 1 0 48668 0 -1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_161_529
timestamp 1644511149
transform 1 0 49772 0 -1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_161_541
timestamp 1644511149
transform 1 0 50876 0 -1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_161_553
timestamp 1644511149
transform 1 0 51980 0 -1 90304
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_161_559
timestamp 1644511149
transform 1 0 52532 0 -1 90304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_161_561
timestamp 1644511149
transform 1 0 52716 0 -1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_161_573
timestamp 1644511149
transform 1 0 53820 0 -1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_161_585
timestamp 1644511149
transform 1 0 54924 0 -1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_161_597
timestamp 1644511149
transform 1 0 56028 0 -1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_161_609
timestamp 1644511149
transform 1 0 57132 0 -1 90304
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_161_615
timestamp 1644511149
transform 1 0 57684 0 -1 90304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_161_617
timestamp 1644511149
transform 1 0 57868 0 -1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_161_629
timestamp 1644511149
transform 1 0 58972 0 -1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_161_641
timestamp 1644511149
transform 1 0 60076 0 -1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_161_653
timestamp 1644511149
transform 1 0 61180 0 -1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_161_665
timestamp 1644511149
transform 1 0 62284 0 -1 90304
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_161_671
timestamp 1644511149
transform 1 0 62836 0 -1 90304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_161_673
timestamp 1644511149
transform 1 0 63020 0 -1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_161_685
timestamp 1644511149
transform 1 0 64124 0 -1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_161_697
timestamp 1644511149
transform 1 0 65228 0 -1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_161_709
timestamp 1644511149
transform 1 0 66332 0 -1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_161_721
timestamp 1644511149
transform 1 0 67436 0 -1 90304
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_161_727
timestamp 1644511149
transform 1 0 67988 0 -1 90304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_161_729
timestamp 1644511149
transform 1 0 68172 0 -1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_161_741
timestamp 1644511149
transform 1 0 69276 0 -1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_161_753
timestamp 1644511149
transform 1 0 70380 0 -1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_161_765
timestamp 1644511149
transform 1 0 71484 0 -1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_161_777
timestamp 1644511149
transform 1 0 72588 0 -1 90304
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_161_783
timestamp 1644511149
transform 1 0 73140 0 -1 90304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_161_785
timestamp 1644511149
transform 1 0 73324 0 -1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_161_797
timestamp 1644511149
transform 1 0 74428 0 -1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_161_809
timestamp 1644511149
transform 1 0 75532 0 -1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_161_821
timestamp 1644511149
transform 1 0 76636 0 -1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_161_833
timestamp 1644511149
transform 1 0 77740 0 -1 90304
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_161_839
timestamp 1644511149
transform 1 0 78292 0 -1 90304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_161_841
timestamp 1644511149
transform 1 0 78476 0 -1 90304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_162_3
timestamp 1644511149
transform 1 0 1380 0 1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_162_15
timestamp 1644511149
transform 1 0 2484 0 1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_162_27
timestamp 1644511149
transform 1 0 3588 0 1 90304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_162_29
timestamp 1644511149
transform 1 0 3772 0 1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_162_41
timestamp 1644511149
transform 1 0 4876 0 1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_162_53
timestamp 1644511149
transform 1 0 5980 0 1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_162_65
timestamp 1644511149
transform 1 0 7084 0 1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_162_77
timestamp 1644511149
transform 1 0 8188 0 1 90304
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_162_83
timestamp 1644511149
transform 1 0 8740 0 1 90304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_162_85
timestamp 1644511149
transform 1 0 8924 0 1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_162_97
timestamp 1644511149
transform 1 0 10028 0 1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_162_109
timestamp 1644511149
transform 1 0 11132 0 1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_162_121
timestamp 1644511149
transform 1 0 12236 0 1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_162_133
timestamp 1644511149
transform 1 0 13340 0 1 90304
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_162_139
timestamp 1644511149
transform 1 0 13892 0 1 90304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_162_141
timestamp 1644511149
transform 1 0 14076 0 1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_162_153
timestamp 1644511149
transform 1 0 15180 0 1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_162_165
timestamp 1644511149
transform 1 0 16284 0 1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_162_177
timestamp 1644511149
transform 1 0 17388 0 1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_162_189
timestamp 1644511149
transform 1 0 18492 0 1 90304
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_162_195
timestamp 1644511149
transform 1 0 19044 0 1 90304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_162_197
timestamp 1644511149
transform 1 0 19228 0 1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_162_209
timestamp 1644511149
transform 1 0 20332 0 1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_162_221
timestamp 1644511149
transform 1 0 21436 0 1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_162_233
timestamp 1644511149
transform 1 0 22540 0 1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_162_245
timestamp 1644511149
transform 1 0 23644 0 1 90304
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_162_251
timestamp 1644511149
transform 1 0 24196 0 1 90304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_162_253
timestamp 1644511149
transform 1 0 24380 0 1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_162_265
timestamp 1644511149
transform 1 0 25484 0 1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_162_277
timestamp 1644511149
transform 1 0 26588 0 1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_162_289
timestamp 1644511149
transform 1 0 27692 0 1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_162_301
timestamp 1644511149
transform 1 0 28796 0 1 90304
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_162_307
timestamp 1644511149
transform 1 0 29348 0 1 90304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_162_309
timestamp 1644511149
transform 1 0 29532 0 1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_162_321
timestamp 1644511149
transform 1 0 30636 0 1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_162_333
timestamp 1644511149
transform 1 0 31740 0 1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_162_345
timestamp 1644511149
transform 1 0 32844 0 1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_162_357
timestamp 1644511149
transform 1 0 33948 0 1 90304
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_162_363
timestamp 1644511149
transform 1 0 34500 0 1 90304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_162_365
timestamp 1644511149
transform 1 0 34684 0 1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_162_377
timestamp 1644511149
transform 1 0 35788 0 1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_162_389
timestamp 1644511149
transform 1 0 36892 0 1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_162_401
timestamp 1644511149
transform 1 0 37996 0 1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_162_413
timestamp 1644511149
transform 1 0 39100 0 1 90304
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_162_419
timestamp 1644511149
transform 1 0 39652 0 1 90304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_162_421
timestamp 1644511149
transform 1 0 39836 0 1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_162_433
timestamp 1644511149
transform 1 0 40940 0 1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_162_445
timestamp 1644511149
transform 1 0 42044 0 1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_162_457
timestamp 1644511149
transform 1 0 43148 0 1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_162_469
timestamp 1644511149
transform 1 0 44252 0 1 90304
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_162_475
timestamp 1644511149
transform 1 0 44804 0 1 90304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_162_477
timestamp 1644511149
transform 1 0 44988 0 1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_162_489
timestamp 1644511149
transform 1 0 46092 0 1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_162_501
timestamp 1644511149
transform 1 0 47196 0 1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_162_513
timestamp 1644511149
transform 1 0 48300 0 1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_162_525
timestamp 1644511149
transform 1 0 49404 0 1 90304
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_162_531
timestamp 1644511149
transform 1 0 49956 0 1 90304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_162_533
timestamp 1644511149
transform 1 0 50140 0 1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_162_545
timestamp 1644511149
transform 1 0 51244 0 1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_162_557
timestamp 1644511149
transform 1 0 52348 0 1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_162_569
timestamp 1644511149
transform 1 0 53452 0 1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_162_581
timestamp 1644511149
transform 1 0 54556 0 1 90304
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_162_587
timestamp 1644511149
transform 1 0 55108 0 1 90304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_162_589
timestamp 1644511149
transform 1 0 55292 0 1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_162_601
timestamp 1644511149
transform 1 0 56396 0 1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_162_613
timestamp 1644511149
transform 1 0 57500 0 1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_162_625
timestamp 1644511149
transform 1 0 58604 0 1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_162_637
timestamp 1644511149
transform 1 0 59708 0 1 90304
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_162_643
timestamp 1644511149
transform 1 0 60260 0 1 90304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_162_645
timestamp 1644511149
transform 1 0 60444 0 1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_162_657
timestamp 1644511149
transform 1 0 61548 0 1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_162_669
timestamp 1644511149
transform 1 0 62652 0 1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_162_681
timestamp 1644511149
transform 1 0 63756 0 1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_162_693
timestamp 1644511149
transform 1 0 64860 0 1 90304
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_162_699
timestamp 1644511149
transform 1 0 65412 0 1 90304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_162_701
timestamp 1644511149
transform 1 0 65596 0 1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_162_713
timestamp 1644511149
transform 1 0 66700 0 1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_162_725
timestamp 1644511149
transform 1 0 67804 0 1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_162_737
timestamp 1644511149
transform 1 0 68908 0 1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_162_749
timestamp 1644511149
transform 1 0 70012 0 1 90304
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_162_755
timestamp 1644511149
transform 1 0 70564 0 1 90304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_162_757
timestamp 1644511149
transform 1 0 70748 0 1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_162_769
timestamp 1644511149
transform 1 0 71852 0 1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_162_781
timestamp 1644511149
transform 1 0 72956 0 1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_162_793
timestamp 1644511149
transform 1 0 74060 0 1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_162_805
timestamp 1644511149
transform 1 0 75164 0 1 90304
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_162_811
timestamp 1644511149
transform 1 0 75716 0 1 90304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_162_813
timestamp 1644511149
transform 1 0 75900 0 1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_162_825
timestamp 1644511149
transform 1 0 77004 0 1 90304
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_162_833
timestamp 1644511149
transform 1 0 77740 0 1 90304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_162_838
timestamp 1644511149
transform 1 0 78200 0 1 90304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_163_3
timestamp 1644511149
transform 1 0 1380 0 -1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_163_15
timestamp 1644511149
transform 1 0 2484 0 -1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_163_27
timestamp 1644511149
transform 1 0 3588 0 -1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_163_39
timestamp 1644511149
transform 1 0 4692 0 -1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_163_51
timestamp 1644511149
transform 1 0 5796 0 -1 91392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_163_55
timestamp 1644511149
transform 1 0 6164 0 -1 91392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_163_57
timestamp 1644511149
transform 1 0 6348 0 -1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_163_69
timestamp 1644511149
transform 1 0 7452 0 -1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_163_81
timestamp 1644511149
transform 1 0 8556 0 -1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_163_93
timestamp 1644511149
transform 1 0 9660 0 -1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_163_105
timestamp 1644511149
transform 1 0 10764 0 -1 91392
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_163_111
timestamp 1644511149
transform 1 0 11316 0 -1 91392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_163_113
timestamp 1644511149
transform 1 0 11500 0 -1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_163_125
timestamp 1644511149
transform 1 0 12604 0 -1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_163_137
timestamp 1644511149
transform 1 0 13708 0 -1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_163_149
timestamp 1644511149
transform 1 0 14812 0 -1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_163_161
timestamp 1644511149
transform 1 0 15916 0 -1 91392
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_163_167
timestamp 1644511149
transform 1 0 16468 0 -1 91392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_163_169
timestamp 1644511149
transform 1 0 16652 0 -1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_163_181
timestamp 1644511149
transform 1 0 17756 0 -1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_163_193
timestamp 1644511149
transform 1 0 18860 0 -1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_163_205
timestamp 1644511149
transform 1 0 19964 0 -1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_163_217
timestamp 1644511149
transform 1 0 21068 0 -1 91392
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_163_223
timestamp 1644511149
transform 1 0 21620 0 -1 91392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_163_225
timestamp 1644511149
transform 1 0 21804 0 -1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_163_237
timestamp 1644511149
transform 1 0 22908 0 -1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_163_249
timestamp 1644511149
transform 1 0 24012 0 -1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_163_261
timestamp 1644511149
transform 1 0 25116 0 -1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_163_273
timestamp 1644511149
transform 1 0 26220 0 -1 91392
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_163_279
timestamp 1644511149
transform 1 0 26772 0 -1 91392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_163_281
timestamp 1644511149
transform 1 0 26956 0 -1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_163_293
timestamp 1644511149
transform 1 0 28060 0 -1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_163_305
timestamp 1644511149
transform 1 0 29164 0 -1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_163_317
timestamp 1644511149
transform 1 0 30268 0 -1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_163_329
timestamp 1644511149
transform 1 0 31372 0 -1 91392
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_163_335
timestamp 1644511149
transform 1 0 31924 0 -1 91392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_163_337
timestamp 1644511149
transform 1 0 32108 0 -1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_163_349
timestamp 1644511149
transform 1 0 33212 0 -1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_163_361
timestamp 1644511149
transform 1 0 34316 0 -1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_163_373
timestamp 1644511149
transform 1 0 35420 0 -1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_163_385
timestamp 1644511149
transform 1 0 36524 0 -1 91392
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_163_391
timestamp 1644511149
transform 1 0 37076 0 -1 91392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_163_393
timestamp 1644511149
transform 1 0 37260 0 -1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_163_405
timestamp 1644511149
transform 1 0 38364 0 -1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_163_417
timestamp 1644511149
transform 1 0 39468 0 -1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_163_429
timestamp 1644511149
transform 1 0 40572 0 -1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_163_441
timestamp 1644511149
transform 1 0 41676 0 -1 91392
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_163_447
timestamp 1644511149
transform 1 0 42228 0 -1 91392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_163_449
timestamp 1644511149
transform 1 0 42412 0 -1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_163_461
timestamp 1644511149
transform 1 0 43516 0 -1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_163_473
timestamp 1644511149
transform 1 0 44620 0 -1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_163_485
timestamp 1644511149
transform 1 0 45724 0 -1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_163_497
timestamp 1644511149
transform 1 0 46828 0 -1 91392
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_163_503
timestamp 1644511149
transform 1 0 47380 0 -1 91392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_163_505
timestamp 1644511149
transform 1 0 47564 0 -1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_163_517
timestamp 1644511149
transform 1 0 48668 0 -1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_163_529
timestamp 1644511149
transform 1 0 49772 0 -1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_163_541
timestamp 1644511149
transform 1 0 50876 0 -1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_163_553
timestamp 1644511149
transform 1 0 51980 0 -1 91392
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_163_559
timestamp 1644511149
transform 1 0 52532 0 -1 91392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_163_561
timestamp 1644511149
transform 1 0 52716 0 -1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_163_573
timestamp 1644511149
transform 1 0 53820 0 -1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_163_585
timestamp 1644511149
transform 1 0 54924 0 -1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_163_597
timestamp 1644511149
transform 1 0 56028 0 -1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_163_609
timestamp 1644511149
transform 1 0 57132 0 -1 91392
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_163_615
timestamp 1644511149
transform 1 0 57684 0 -1 91392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_163_617
timestamp 1644511149
transform 1 0 57868 0 -1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_163_629
timestamp 1644511149
transform 1 0 58972 0 -1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_163_641
timestamp 1644511149
transform 1 0 60076 0 -1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_163_653
timestamp 1644511149
transform 1 0 61180 0 -1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_163_665
timestamp 1644511149
transform 1 0 62284 0 -1 91392
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_163_671
timestamp 1644511149
transform 1 0 62836 0 -1 91392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_163_673
timestamp 1644511149
transform 1 0 63020 0 -1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_163_685
timestamp 1644511149
transform 1 0 64124 0 -1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_163_697
timestamp 1644511149
transform 1 0 65228 0 -1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_163_709
timestamp 1644511149
transform 1 0 66332 0 -1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_163_721
timestamp 1644511149
transform 1 0 67436 0 -1 91392
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_163_727
timestamp 1644511149
transform 1 0 67988 0 -1 91392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_163_729
timestamp 1644511149
transform 1 0 68172 0 -1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_163_741
timestamp 1644511149
transform 1 0 69276 0 -1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_163_753
timestamp 1644511149
transform 1 0 70380 0 -1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_163_765
timestamp 1644511149
transform 1 0 71484 0 -1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_163_777
timestamp 1644511149
transform 1 0 72588 0 -1 91392
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_163_783
timestamp 1644511149
transform 1 0 73140 0 -1 91392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_163_785
timestamp 1644511149
transform 1 0 73324 0 -1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_163_797
timestamp 1644511149
transform 1 0 74428 0 -1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_163_809
timestamp 1644511149
transform 1 0 75532 0 -1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_163_821
timestamp 1644511149
transform 1 0 76636 0 -1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_163_833
timestamp 1644511149
transform 1 0 77740 0 -1 91392
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_163_839
timestamp 1644511149
transform 1 0 78292 0 -1 91392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_163_841
timestamp 1644511149
transform 1 0 78476 0 -1 91392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_164_3
timestamp 1644511149
transform 1 0 1380 0 1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_164_15
timestamp 1644511149
transform 1 0 2484 0 1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_164_27
timestamp 1644511149
transform 1 0 3588 0 1 91392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_164_29
timestamp 1644511149
transform 1 0 3772 0 1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_164_41
timestamp 1644511149
transform 1 0 4876 0 1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_164_53
timestamp 1644511149
transform 1 0 5980 0 1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_164_65
timestamp 1644511149
transform 1 0 7084 0 1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_164_77
timestamp 1644511149
transform 1 0 8188 0 1 91392
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_164_83
timestamp 1644511149
transform 1 0 8740 0 1 91392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_164_85
timestamp 1644511149
transform 1 0 8924 0 1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_164_97
timestamp 1644511149
transform 1 0 10028 0 1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_164_109
timestamp 1644511149
transform 1 0 11132 0 1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_164_121
timestamp 1644511149
transform 1 0 12236 0 1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_164_133
timestamp 1644511149
transform 1 0 13340 0 1 91392
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_164_139
timestamp 1644511149
transform 1 0 13892 0 1 91392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_164_141
timestamp 1644511149
transform 1 0 14076 0 1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_164_153
timestamp 1644511149
transform 1 0 15180 0 1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_164_165
timestamp 1644511149
transform 1 0 16284 0 1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_164_177
timestamp 1644511149
transform 1 0 17388 0 1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_164_189
timestamp 1644511149
transform 1 0 18492 0 1 91392
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_164_195
timestamp 1644511149
transform 1 0 19044 0 1 91392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_164_197
timestamp 1644511149
transform 1 0 19228 0 1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_164_209
timestamp 1644511149
transform 1 0 20332 0 1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_164_221
timestamp 1644511149
transform 1 0 21436 0 1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_164_233
timestamp 1644511149
transform 1 0 22540 0 1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_164_245
timestamp 1644511149
transform 1 0 23644 0 1 91392
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_164_251
timestamp 1644511149
transform 1 0 24196 0 1 91392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_164_253
timestamp 1644511149
transform 1 0 24380 0 1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_164_265
timestamp 1644511149
transform 1 0 25484 0 1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_164_277
timestamp 1644511149
transform 1 0 26588 0 1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_164_289
timestamp 1644511149
transform 1 0 27692 0 1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_164_301
timestamp 1644511149
transform 1 0 28796 0 1 91392
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_164_307
timestamp 1644511149
transform 1 0 29348 0 1 91392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_164_309
timestamp 1644511149
transform 1 0 29532 0 1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_164_321
timestamp 1644511149
transform 1 0 30636 0 1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_164_333
timestamp 1644511149
transform 1 0 31740 0 1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_164_345
timestamp 1644511149
transform 1 0 32844 0 1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_164_357
timestamp 1644511149
transform 1 0 33948 0 1 91392
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_164_363
timestamp 1644511149
transform 1 0 34500 0 1 91392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_164_365
timestamp 1644511149
transform 1 0 34684 0 1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_164_377
timestamp 1644511149
transform 1 0 35788 0 1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_164_389
timestamp 1644511149
transform 1 0 36892 0 1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_164_401
timestamp 1644511149
transform 1 0 37996 0 1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_164_413
timestamp 1644511149
transform 1 0 39100 0 1 91392
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_164_419
timestamp 1644511149
transform 1 0 39652 0 1 91392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_164_421
timestamp 1644511149
transform 1 0 39836 0 1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_164_433
timestamp 1644511149
transform 1 0 40940 0 1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_164_445
timestamp 1644511149
transform 1 0 42044 0 1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_164_457
timestamp 1644511149
transform 1 0 43148 0 1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_164_469
timestamp 1644511149
transform 1 0 44252 0 1 91392
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_164_475
timestamp 1644511149
transform 1 0 44804 0 1 91392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_164_477
timestamp 1644511149
transform 1 0 44988 0 1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_164_489
timestamp 1644511149
transform 1 0 46092 0 1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_164_501
timestamp 1644511149
transform 1 0 47196 0 1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_164_513
timestamp 1644511149
transform 1 0 48300 0 1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_164_525
timestamp 1644511149
transform 1 0 49404 0 1 91392
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_164_531
timestamp 1644511149
transform 1 0 49956 0 1 91392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_164_533
timestamp 1644511149
transform 1 0 50140 0 1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_164_545
timestamp 1644511149
transform 1 0 51244 0 1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_164_557
timestamp 1644511149
transform 1 0 52348 0 1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_164_569
timestamp 1644511149
transform 1 0 53452 0 1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_164_581
timestamp 1644511149
transform 1 0 54556 0 1 91392
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_164_587
timestamp 1644511149
transform 1 0 55108 0 1 91392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_164_589
timestamp 1644511149
transform 1 0 55292 0 1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_164_601
timestamp 1644511149
transform 1 0 56396 0 1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_164_613
timestamp 1644511149
transform 1 0 57500 0 1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_164_625
timestamp 1644511149
transform 1 0 58604 0 1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_164_637
timestamp 1644511149
transform 1 0 59708 0 1 91392
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_164_643
timestamp 1644511149
transform 1 0 60260 0 1 91392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_164_645
timestamp 1644511149
transform 1 0 60444 0 1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_164_657
timestamp 1644511149
transform 1 0 61548 0 1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_164_669
timestamp 1644511149
transform 1 0 62652 0 1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_164_681
timestamp 1644511149
transform 1 0 63756 0 1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_164_693
timestamp 1644511149
transform 1 0 64860 0 1 91392
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_164_699
timestamp 1644511149
transform 1 0 65412 0 1 91392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_164_701
timestamp 1644511149
transform 1 0 65596 0 1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_164_713
timestamp 1644511149
transform 1 0 66700 0 1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_164_725
timestamp 1644511149
transform 1 0 67804 0 1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_164_737
timestamp 1644511149
transform 1 0 68908 0 1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_164_749
timestamp 1644511149
transform 1 0 70012 0 1 91392
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_164_755
timestamp 1644511149
transform 1 0 70564 0 1 91392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_164_757
timestamp 1644511149
transform 1 0 70748 0 1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_164_769
timestamp 1644511149
transform 1 0 71852 0 1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_164_781
timestamp 1644511149
transform 1 0 72956 0 1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_164_793
timestamp 1644511149
transform 1 0 74060 0 1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_164_805
timestamp 1644511149
transform 1 0 75164 0 1 91392
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_164_811
timestamp 1644511149
transform 1 0 75716 0 1 91392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_164_813
timestamp 1644511149
transform 1 0 75900 0 1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_164_825
timestamp 1644511149
transform 1 0 77004 0 1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_164_837
timestamp 1644511149
transform 1 0 78108 0 1 91392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_164_841
timestamp 1644511149
transform 1 0 78476 0 1 91392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_165_3
timestamp 1644511149
transform 1 0 1380 0 -1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_165_15
timestamp 1644511149
transform 1 0 2484 0 -1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_165_27
timestamp 1644511149
transform 1 0 3588 0 -1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_165_39
timestamp 1644511149
transform 1 0 4692 0 -1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_165_51
timestamp 1644511149
transform 1 0 5796 0 -1 92480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_165_55
timestamp 1644511149
transform 1 0 6164 0 -1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_165_57
timestamp 1644511149
transform 1 0 6348 0 -1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_165_69
timestamp 1644511149
transform 1 0 7452 0 -1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_165_81
timestamp 1644511149
transform 1 0 8556 0 -1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_165_93
timestamp 1644511149
transform 1 0 9660 0 -1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_165_105
timestamp 1644511149
transform 1 0 10764 0 -1 92480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_165_111
timestamp 1644511149
transform 1 0 11316 0 -1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_165_113
timestamp 1644511149
transform 1 0 11500 0 -1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_165_125
timestamp 1644511149
transform 1 0 12604 0 -1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_165_137
timestamp 1644511149
transform 1 0 13708 0 -1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_165_149
timestamp 1644511149
transform 1 0 14812 0 -1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_165_161
timestamp 1644511149
transform 1 0 15916 0 -1 92480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_165_167
timestamp 1644511149
transform 1 0 16468 0 -1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_165_169
timestamp 1644511149
transform 1 0 16652 0 -1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_165_181
timestamp 1644511149
transform 1 0 17756 0 -1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_165_193
timestamp 1644511149
transform 1 0 18860 0 -1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_165_205
timestamp 1644511149
transform 1 0 19964 0 -1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_165_217
timestamp 1644511149
transform 1 0 21068 0 -1 92480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_165_223
timestamp 1644511149
transform 1 0 21620 0 -1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_165_225
timestamp 1644511149
transform 1 0 21804 0 -1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_165_237
timestamp 1644511149
transform 1 0 22908 0 -1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_165_249
timestamp 1644511149
transform 1 0 24012 0 -1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_165_261
timestamp 1644511149
transform 1 0 25116 0 -1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_165_273
timestamp 1644511149
transform 1 0 26220 0 -1 92480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_165_279
timestamp 1644511149
transform 1 0 26772 0 -1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_165_281
timestamp 1644511149
transform 1 0 26956 0 -1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_165_293
timestamp 1644511149
transform 1 0 28060 0 -1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_165_305
timestamp 1644511149
transform 1 0 29164 0 -1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_165_317
timestamp 1644511149
transform 1 0 30268 0 -1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_165_329
timestamp 1644511149
transform 1 0 31372 0 -1 92480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_165_335
timestamp 1644511149
transform 1 0 31924 0 -1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_165_337
timestamp 1644511149
transform 1 0 32108 0 -1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_165_349
timestamp 1644511149
transform 1 0 33212 0 -1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_165_361
timestamp 1644511149
transform 1 0 34316 0 -1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_165_373
timestamp 1644511149
transform 1 0 35420 0 -1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_165_385
timestamp 1644511149
transform 1 0 36524 0 -1 92480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_165_391
timestamp 1644511149
transform 1 0 37076 0 -1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_165_393
timestamp 1644511149
transform 1 0 37260 0 -1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_165_405
timestamp 1644511149
transform 1 0 38364 0 -1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_165_417
timestamp 1644511149
transform 1 0 39468 0 -1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_165_429
timestamp 1644511149
transform 1 0 40572 0 -1 92480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_165_440
timestamp 1644511149
transform 1 0 41584 0 -1 92480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_165_449
timestamp 1644511149
transform 1 0 42412 0 -1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_165_461
timestamp 1644511149
transform 1 0 43516 0 -1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_165_473
timestamp 1644511149
transform 1 0 44620 0 -1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_165_485
timestamp 1644511149
transform 1 0 45724 0 -1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_165_497
timestamp 1644511149
transform 1 0 46828 0 -1 92480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_165_503
timestamp 1644511149
transform 1 0 47380 0 -1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_165_505
timestamp 1644511149
transform 1 0 47564 0 -1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_165_517
timestamp 1644511149
transform 1 0 48668 0 -1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_165_529
timestamp 1644511149
transform 1 0 49772 0 -1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_165_541
timestamp 1644511149
transform 1 0 50876 0 -1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_165_553
timestamp 1644511149
transform 1 0 51980 0 -1 92480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_165_559
timestamp 1644511149
transform 1 0 52532 0 -1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_165_561
timestamp 1644511149
transform 1 0 52716 0 -1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_165_573
timestamp 1644511149
transform 1 0 53820 0 -1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_165_585
timestamp 1644511149
transform 1 0 54924 0 -1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_165_597
timestamp 1644511149
transform 1 0 56028 0 -1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_165_609
timestamp 1644511149
transform 1 0 57132 0 -1 92480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_165_615
timestamp 1644511149
transform 1 0 57684 0 -1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_165_617
timestamp 1644511149
transform 1 0 57868 0 -1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_165_629
timestamp 1644511149
transform 1 0 58972 0 -1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_165_641
timestamp 1644511149
transform 1 0 60076 0 -1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_165_653
timestamp 1644511149
transform 1 0 61180 0 -1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_165_665
timestamp 1644511149
transform 1 0 62284 0 -1 92480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_165_671
timestamp 1644511149
transform 1 0 62836 0 -1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_165_673
timestamp 1644511149
transform 1 0 63020 0 -1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_165_685
timestamp 1644511149
transform 1 0 64124 0 -1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_165_697
timestamp 1644511149
transform 1 0 65228 0 -1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_165_709
timestamp 1644511149
transform 1 0 66332 0 -1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_165_721
timestamp 1644511149
transform 1 0 67436 0 -1 92480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_165_727
timestamp 1644511149
transform 1 0 67988 0 -1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_165_729
timestamp 1644511149
transform 1 0 68172 0 -1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_165_741
timestamp 1644511149
transform 1 0 69276 0 -1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_165_753
timestamp 1644511149
transform 1 0 70380 0 -1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_165_765
timestamp 1644511149
transform 1 0 71484 0 -1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_165_777
timestamp 1644511149
transform 1 0 72588 0 -1 92480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_165_783
timestamp 1644511149
transform 1 0 73140 0 -1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_165_785
timestamp 1644511149
transform 1 0 73324 0 -1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_165_797
timestamp 1644511149
transform 1 0 74428 0 -1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_165_809
timestamp 1644511149
transform 1 0 75532 0 -1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_165_821
timestamp 1644511149
transform 1 0 76636 0 -1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_165_833
timestamp 1644511149
transform 1 0 77740 0 -1 92480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_165_839
timestamp 1644511149
transform 1 0 78292 0 -1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_165_841
timestamp 1644511149
transform 1 0 78476 0 -1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_166_3
timestamp 1644511149
transform 1 0 1380 0 1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_166_15
timestamp 1644511149
transform 1 0 2484 0 1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_166_27
timestamp 1644511149
transform 1 0 3588 0 1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_166_29
timestamp 1644511149
transform 1 0 3772 0 1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_166_41
timestamp 1644511149
transform 1 0 4876 0 1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_166_53
timestamp 1644511149
transform 1 0 5980 0 1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_166_65
timestamp 1644511149
transform 1 0 7084 0 1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_166_77
timestamp 1644511149
transform 1 0 8188 0 1 92480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_166_83
timestamp 1644511149
transform 1 0 8740 0 1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_166_85
timestamp 1644511149
transform 1 0 8924 0 1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_166_97
timestamp 1644511149
transform 1 0 10028 0 1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_166_109
timestamp 1644511149
transform 1 0 11132 0 1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_166_121
timestamp 1644511149
transform 1 0 12236 0 1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_166_133
timestamp 1644511149
transform 1 0 13340 0 1 92480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_166_139
timestamp 1644511149
transform 1 0 13892 0 1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_166_141
timestamp 1644511149
transform 1 0 14076 0 1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_166_153
timestamp 1644511149
transform 1 0 15180 0 1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_166_165
timestamp 1644511149
transform 1 0 16284 0 1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_166_177
timestamp 1644511149
transform 1 0 17388 0 1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_166_189
timestamp 1644511149
transform 1 0 18492 0 1 92480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_166_195
timestamp 1644511149
transform 1 0 19044 0 1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_166_197
timestamp 1644511149
transform 1 0 19228 0 1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_166_209
timestamp 1644511149
transform 1 0 20332 0 1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_166_221
timestamp 1644511149
transform 1 0 21436 0 1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_166_233
timestamp 1644511149
transform 1 0 22540 0 1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_166_245
timestamp 1644511149
transform 1 0 23644 0 1 92480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_166_251
timestamp 1644511149
transform 1 0 24196 0 1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_166_253
timestamp 1644511149
transform 1 0 24380 0 1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_166_265
timestamp 1644511149
transform 1 0 25484 0 1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_166_277
timestamp 1644511149
transform 1 0 26588 0 1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_166_289
timestamp 1644511149
transform 1 0 27692 0 1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_166_301
timestamp 1644511149
transform 1 0 28796 0 1 92480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_166_307
timestamp 1644511149
transform 1 0 29348 0 1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_166_309
timestamp 1644511149
transform 1 0 29532 0 1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_166_321
timestamp 1644511149
transform 1 0 30636 0 1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_166_333
timestamp 1644511149
transform 1 0 31740 0 1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_166_345
timestamp 1644511149
transform 1 0 32844 0 1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_166_357
timestamp 1644511149
transform 1 0 33948 0 1 92480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_166_363
timestamp 1644511149
transform 1 0 34500 0 1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_166_365
timestamp 1644511149
transform 1 0 34684 0 1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_166_377
timestamp 1644511149
transform 1 0 35788 0 1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_166_389
timestamp 1644511149
transform 1 0 36892 0 1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_166_401
timestamp 1644511149
transform 1 0 37996 0 1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_166_413
timestamp 1644511149
transform 1 0 39100 0 1 92480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_166_419
timestamp 1644511149
transform 1 0 39652 0 1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_166_421
timestamp 1644511149
transform 1 0 39836 0 1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_166_433
timestamp 1644511149
transform 1 0 40940 0 1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_166_445
timestamp 1644511149
transform 1 0 42044 0 1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_166_457
timestamp 1644511149
transform 1 0 43148 0 1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_166_469
timestamp 1644511149
transform 1 0 44252 0 1 92480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_166_475
timestamp 1644511149
transform 1 0 44804 0 1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_166_477
timestamp 1644511149
transform 1 0 44988 0 1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_166_489
timestamp 1644511149
transform 1 0 46092 0 1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_166_501
timestamp 1644511149
transform 1 0 47196 0 1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_166_513
timestamp 1644511149
transform 1 0 48300 0 1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_166_525
timestamp 1644511149
transform 1 0 49404 0 1 92480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_166_531
timestamp 1644511149
transform 1 0 49956 0 1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_166_533
timestamp 1644511149
transform 1 0 50140 0 1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_166_545
timestamp 1644511149
transform 1 0 51244 0 1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_166_557
timestamp 1644511149
transform 1 0 52348 0 1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_166_569
timestamp 1644511149
transform 1 0 53452 0 1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_166_581
timestamp 1644511149
transform 1 0 54556 0 1 92480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_166_587
timestamp 1644511149
transform 1 0 55108 0 1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_166_589
timestamp 1644511149
transform 1 0 55292 0 1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_166_601
timestamp 1644511149
transform 1 0 56396 0 1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_166_613
timestamp 1644511149
transform 1 0 57500 0 1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_166_625
timestamp 1644511149
transform 1 0 58604 0 1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_166_637
timestamp 1644511149
transform 1 0 59708 0 1 92480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_166_643
timestamp 1644511149
transform 1 0 60260 0 1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_166_645
timestamp 1644511149
transform 1 0 60444 0 1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_166_657
timestamp 1644511149
transform 1 0 61548 0 1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_166_669
timestamp 1644511149
transform 1 0 62652 0 1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_166_681
timestamp 1644511149
transform 1 0 63756 0 1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_166_693
timestamp 1644511149
transform 1 0 64860 0 1 92480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_166_699
timestamp 1644511149
transform 1 0 65412 0 1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_166_701
timestamp 1644511149
transform 1 0 65596 0 1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_166_713
timestamp 1644511149
transform 1 0 66700 0 1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_166_725
timestamp 1644511149
transform 1 0 67804 0 1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_166_737
timestamp 1644511149
transform 1 0 68908 0 1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_166_749
timestamp 1644511149
transform 1 0 70012 0 1 92480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_166_755
timestamp 1644511149
transform 1 0 70564 0 1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_166_757
timestamp 1644511149
transform 1 0 70748 0 1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_166_769
timestamp 1644511149
transform 1 0 71852 0 1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_166_781
timestamp 1644511149
transform 1 0 72956 0 1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_166_793
timestamp 1644511149
transform 1 0 74060 0 1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_166_805
timestamp 1644511149
transform 1 0 75164 0 1 92480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_166_811
timestamp 1644511149
transform 1 0 75716 0 1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_166_813
timestamp 1644511149
transform 1 0 75900 0 1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_166_825
timestamp 1644511149
transform 1 0 77004 0 1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_166_837
timestamp 1644511149
transform 1 0 78108 0 1 92480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_166_841
timestamp 1644511149
transform 1 0 78476 0 1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_167_3
timestamp 1644511149
transform 1 0 1380 0 -1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_167_15
timestamp 1644511149
transform 1 0 2484 0 -1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_167_27
timestamp 1644511149
transform 1 0 3588 0 -1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_167_39
timestamp 1644511149
transform 1 0 4692 0 -1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_167_51
timestamp 1644511149
transform 1 0 5796 0 -1 93568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_167_55
timestamp 1644511149
transform 1 0 6164 0 -1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_167_57
timestamp 1644511149
transform 1 0 6348 0 -1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_167_69
timestamp 1644511149
transform 1 0 7452 0 -1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_167_81
timestamp 1644511149
transform 1 0 8556 0 -1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_167_93
timestamp 1644511149
transform 1 0 9660 0 -1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_167_105
timestamp 1644511149
transform 1 0 10764 0 -1 93568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_167_111
timestamp 1644511149
transform 1 0 11316 0 -1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_167_113
timestamp 1644511149
transform 1 0 11500 0 -1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_167_125
timestamp 1644511149
transform 1 0 12604 0 -1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_167_137
timestamp 1644511149
transform 1 0 13708 0 -1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_167_149
timestamp 1644511149
transform 1 0 14812 0 -1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_167_161
timestamp 1644511149
transform 1 0 15916 0 -1 93568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_167_167
timestamp 1644511149
transform 1 0 16468 0 -1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_167_169
timestamp 1644511149
transform 1 0 16652 0 -1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_167_181
timestamp 1644511149
transform 1 0 17756 0 -1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_167_193
timestamp 1644511149
transform 1 0 18860 0 -1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_167_205
timestamp 1644511149
transform 1 0 19964 0 -1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_167_217
timestamp 1644511149
transform 1 0 21068 0 -1 93568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_167_223
timestamp 1644511149
transform 1 0 21620 0 -1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_167_225
timestamp 1644511149
transform 1 0 21804 0 -1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_167_237
timestamp 1644511149
transform 1 0 22908 0 -1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_167_249
timestamp 1644511149
transform 1 0 24012 0 -1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_167_261
timestamp 1644511149
transform 1 0 25116 0 -1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_167_273
timestamp 1644511149
transform 1 0 26220 0 -1 93568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_167_279
timestamp 1644511149
transform 1 0 26772 0 -1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_167_281
timestamp 1644511149
transform 1 0 26956 0 -1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_167_293
timestamp 1644511149
transform 1 0 28060 0 -1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_167_305
timestamp 1644511149
transform 1 0 29164 0 -1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_167_317
timestamp 1644511149
transform 1 0 30268 0 -1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_167_329
timestamp 1644511149
transform 1 0 31372 0 -1 93568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_167_335
timestamp 1644511149
transform 1 0 31924 0 -1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_167_337
timestamp 1644511149
transform 1 0 32108 0 -1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_167_349
timestamp 1644511149
transform 1 0 33212 0 -1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_167_361
timestamp 1644511149
transform 1 0 34316 0 -1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_167_373
timestamp 1644511149
transform 1 0 35420 0 -1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_167_385
timestamp 1644511149
transform 1 0 36524 0 -1 93568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_167_391
timestamp 1644511149
transform 1 0 37076 0 -1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_167_393
timestamp 1644511149
transform 1 0 37260 0 -1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_167_405
timestamp 1644511149
transform 1 0 38364 0 -1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_167_417
timestamp 1644511149
transform 1 0 39468 0 -1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_167_429
timestamp 1644511149
transform 1 0 40572 0 -1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_167_441
timestamp 1644511149
transform 1 0 41676 0 -1 93568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_167_447
timestamp 1644511149
transform 1 0 42228 0 -1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_167_449
timestamp 1644511149
transform 1 0 42412 0 -1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_167_461
timestamp 1644511149
transform 1 0 43516 0 -1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_167_473
timestamp 1644511149
transform 1 0 44620 0 -1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_167_485
timestamp 1644511149
transform 1 0 45724 0 -1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_167_497
timestamp 1644511149
transform 1 0 46828 0 -1 93568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_167_503
timestamp 1644511149
transform 1 0 47380 0 -1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_167_505
timestamp 1644511149
transform 1 0 47564 0 -1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_167_517
timestamp 1644511149
transform 1 0 48668 0 -1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_167_529
timestamp 1644511149
transform 1 0 49772 0 -1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_167_541
timestamp 1644511149
transform 1 0 50876 0 -1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_167_553
timestamp 1644511149
transform 1 0 51980 0 -1 93568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_167_559
timestamp 1644511149
transform 1 0 52532 0 -1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_167_561
timestamp 1644511149
transform 1 0 52716 0 -1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_167_573
timestamp 1644511149
transform 1 0 53820 0 -1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_167_585
timestamp 1644511149
transform 1 0 54924 0 -1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_167_597
timestamp 1644511149
transform 1 0 56028 0 -1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_167_609
timestamp 1644511149
transform 1 0 57132 0 -1 93568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_167_615
timestamp 1644511149
transform 1 0 57684 0 -1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_167_617
timestamp 1644511149
transform 1 0 57868 0 -1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_167_629
timestamp 1644511149
transform 1 0 58972 0 -1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_167_641
timestamp 1644511149
transform 1 0 60076 0 -1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_167_653
timestamp 1644511149
transform 1 0 61180 0 -1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_167_665
timestamp 1644511149
transform 1 0 62284 0 -1 93568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_167_671
timestamp 1644511149
transform 1 0 62836 0 -1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_167_673
timestamp 1644511149
transform 1 0 63020 0 -1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_167_685
timestamp 1644511149
transform 1 0 64124 0 -1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_167_697
timestamp 1644511149
transform 1 0 65228 0 -1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_167_709
timestamp 1644511149
transform 1 0 66332 0 -1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_167_721
timestamp 1644511149
transform 1 0 67436 0 -1 93568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_167_727
timestamp 1644511149
transform 1 0 67988 0 -1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_167_729
timestamp 1644511149
transform 1 0 68172 0 -1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_167_741
timestamp 1644511149
transform 1 0 69276 0 -1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_167_753
timestamp 1644511149
transform 1 0 70380 0 -1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_167_765
timestamp 1644511149
transform 1 0 71484 0 -1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_167_777
timestamp 1644511149
transform 1 0 72588 0 -1 93568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_167_783
timestamp 1644511149
transform 1 0 73140 0 -1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_167_785
timestamp 1644511149
transform 1 0 73324 0 -1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_167_797
timestamp 1644511149
transform 1 0 74428 0 -1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_167_809
timestamp 1644511149
transform 1 0 75532 0 -1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_167_821
timestamp 1644511149
transform 1 0 76636 0 -1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_167_833
timestamp 1644511149
transform 1 0 77740 0 -1 93568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_167_839
timestamp 1644511149
transform 1 0 78292 0 -1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_167_841
timestamp 1644511149
transform 1 0 78476 0 -1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_168_3
timestamp 1644511149
transform 1 0 1380 0 1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_168_15
timestamp 1644511149
transform 1 0 2484 0 1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_168_27
timestamp 1644511149
transform 1 0 3588 0 1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_168_29
timestamp 1644511149
transform 1 0 3772 0 1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_168_41
timestamp 1644511149
transform 1 0 4876 0 1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_168_53
timestamp 1644511149
transform 1 0 5980 0 1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_168_65
timestamp 1644511149
transform 1 0 7084 0 1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_168_77
timestamp 1644511149
transform 1 0 8188 0 1 93568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_168_83
timestamp 1644511149
transform 1 0 8740 0 1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_168_85
timestamp 1644511149
transform 1 0 8924 0 1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_168_97
timestamp 1644511149
transform 1 0 10028 0 1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_168_109
timestamp 1644511149
transform 1 0 11132 0 1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_168_121
timestamp 1644511149
transform 1 0 12236 0 1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_168_133
timestamp 1644511149
transform 1 0 13340 0 1 93568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_168_139
timestamp 1644511149
transform 1 0 13892 0 1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_168_141
timestamp 1644511149
transform 1 0 14076 0 1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_168_153
timestamp 1644511149
transform 1 0 15180 0 1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_168_165
timestamp 1644511149
transform 1 0 16284 0 1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_168_177
timestamp 1644511149
transform 1 0 17388 0 1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_168_189
timestamp 1644511149
transform 1 0 18492 0 1 93568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_168_195
timestamp 1644511149
transform 1 0 19044 0 1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_168_197
timestamp 1644511149
transform 1 0 19228 0 1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_168_209
timestamp 1644511149
transform 1 0 20332 0 1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_168_221
timestamp 1644511149
transform 1 0 21436 0 1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_168_233
timestamp 1644511149
transform 1 0 22540 0 1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_168_245
timestamp 1644511149
transform 1 0 23644 0 1 93568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_168_251
timestamp 1644511149
transform 1 0 24196 0 1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_168_253
timestamp 1644511149
transform 1 0 24380 0 1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_168_265
timestamp 1644511149
transform 1 0 25484 0 1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_168_277
timestamp 1644511149
transform 1 0 26588 0 1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_168_289
timestamp 1644511149
transform 1 0 27692 0 1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_168_301
timestamp 1644511149
transform 1 0 28796 0 1 93568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_168_307
timestamp 1644511149
transform 1 0 29348 0 1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_168_309
timestamp 1644511149
transform 1 0 29532 0 1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_168_321
timestamp 1644511149
transform 1 0 30636 0 1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_168_333
timestamp 1644511149
transform 1 0 31740 0 1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_168_345
timestamp 1644511149
transform 1 0 32844 0 1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_168_357
timestamp 1644511149
transform 1 0 33948 0 1 93568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_168_363
timestamp 1644511149
transform 1 0 34500 0 1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_168_365
timestamp 1644511149
transform 1 0 34684 0 1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_168_377
timestamp 1644511149
transform 1 0 35788 0 1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_168_389
timestamp 1644511149
transform 1 0 36892 0 1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_168_401
timestamp 1644511149
transform 1 0 37996 0 1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_168_413
timestamp 1644511149
transform 1 0 39100 0 1 93568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_168_419
timestamp 1644511149
transform 1 0 39652 0 1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_168_421
timestamp 1644511149
transform 1 0 39836 0 1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_168_433
timestamp 1644511149
transform 1 0 40940 0 1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_168_445
timestamp 1644511149
transform 1 0 42044 0 1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_168_457
timestamp 1644511149
transform 1 0 43148 0 1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_168_469
timestamp 1644511149
transform 1 0 44252 0 1 93568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_168_475
timestamp 1644511149
transform 1 0 44804 0 1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_168_477
timestamp 1644511149
transform 1 0 44988 0 1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_168_489
timestamp 1644511149
transform 1 0 46092 0 1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_168_501
timestamp 1644511149
transform 1 0 47196 0 1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_168_513
timestamp 1644511149
transform 1 0 48300 0 1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_168_525
timestamp 1644511149
transform 1 0 49404 0 1 93568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_168_531
timestamp 1644511149
transform 1 0 49956 0 1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_168_533
timestamp 1644511149
transform 1 0 50140 0 1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_168_545
timestamp 1644511149
transform 1 0 51244 0 1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_168_557
timestamp 1644511149
transform 1 0 52348 0 1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_168_569
timestamp 1644511149
transform 1 0 53452 0 1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_168_581
timestamp 1644511149
transform 1 0 54556 0 1 93568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_168_587
timestamp 1644511149
transform 1 0 55108 0 1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_168_589
timestamp 1644511149
transform 1 0 55292 0 1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_168_601
timestamp 1644511149
transform 1 0 56396 0 1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_168_613
timestamp 1644511149
transform 1 0 57500 0 1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_168_625
timestamp 1644511149
transform 1 0 58604 0 1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_168_637
timestamp 1644511149
transform 1 0 59708 0 1 93568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_168_643
timestamp 1644511149
transform 1 0 60260 0 1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_168_645
timestamp 1644511149
transform 1 0 60444 0 1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_168_657
timestamp 1644511149
transform 1 0 61548 0 1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_168_669
timestamp 1644511149
transform 1 0 62652 0 1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_168_681
timestamp 1644511149
transform 1 0 63756 0 1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_168_693
timestamp 1644511149
transform 1 0 64860 0 1 93568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_168_699
timestamp 1644511149
transform 1 0 65412 0 1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_168_701
timestamp 1644511149
transform 1 0 65596 0 1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_168_713
timestamp 1644511149
transform 1 0 66700 0 1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_168_725
timestamp 1644511149
transform 1 0 67804 0 1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_168_737
timestamp 1644511149
transform 1 0 68908 0 1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_168_749
timestamp 1644511149
transform 1 0 70012 0 1 93568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_168_755
timestamp 1644511149
transform 1 0 70564 0 1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_168_757
timestamp 1644511149
transform 1 0 70748 0 1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_168_769
timestamp 1644511149
transform 1 0 71852 0 1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_168_781
timestamp 1644511149
transform 1 0 72956 0 1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_168_793
timestamp 1644511149
transform 1 0 74060 0 1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_168_805
timestamp 1644511149
transform 1 0 75164 0 1 93568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_168_811
timestamp 1644511149
transform 1 0 75716 0 1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_168_813
timestamp 1644511149
transform 1 0 75900 0 1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_168_825
timestamp 1644511149
transform 1 0 77004 0 1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_168_837
timestamp 1644511149
transform 1 0 78108 0 1 93568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_168_841
timestamp 1644511149
transform 1 0 78476 0 1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_169_7
timestamp 1644511149
transform 1 0 1748 0 -1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_169_19
timestamp 1644511149
transform 1 0 2852 0 -1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_169_31
timestamp 1644511149
transform 1 0 3956 0 -1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_169_43
timestamp 1644511149
transform 1 0 5060 0 -1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_169_55
timestamp 1644511149
transform 1 0 6164 0 -1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_169_57
timestamp 1644511149
transform 1 0 6348 0 -1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_169_69
timestamp 1644511149
transform 1 0 7452 0 -1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_169_81
timestamp 1644511149
transform 1 0 8556 0 -1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_169_93
timestamp 1644511149
transform 1 0 9660 0 -1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_169_105
timestamp 1644511149
transform 1 0 10764 0 -1 94656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_169_111
timestamp 1644511149
transform 1 0 11316 0 -1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_169_113
timestamp 1644511149
transform 1 0 11500 0 -1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_169_125
timestamp 1644511149
transform 1 0 12604 0 -1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_169_137
timestamp 1644511149
transform 1 0 13708 0 -1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_169_149
timestamp 1644511149
transform 1 0 14812 0 -1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_169_161
timestamp 1644511149
transform 1 0 15916 0 -1 94656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_169_167
timestamp 1644511149
transform 1 0 16468 0 -1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_169_169
timestamp 1644511149
transform 1 0 16652 0 -1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_169_181
timestamp 1644511149
transform 1 0 17756 0 -1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_169_193
timestamp 1644511149
transform 1 0 18860 0 -1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_169_205
timestamp 1644511149
transform 1 0 19964 0 -1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_169_217
timestamp 1644511149
transform 1 0 21068 0 -1 94656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_169_223
timestamp 1644511149
transform 1 0 21620 0 -1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_169_225
timestamp 1644511149
transform 1 0 21804 0 -1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_169_237
timestamp 1644511149
transform 1 0 22908 0 -1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_169_249
timestamp 1644511149
transform 1 0 24012 0 -1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_169_261
timestamp 1644511149
transform 1 0 25116 0 -1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_169_273
timestamp 1644511149
transform 1 0 26220 0 -1 94656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_169_279
timestamp 1644511149
transform 1 0 26772 0 -1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_169_281
timestamp 1644511149
transform 1 0 26956 0 -1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_169_293
timestamp 1644511149
transform 1 0 28060 0 -1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_169_305
timestamp 1644511149
transform 1 0 29164 0 -1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_169_317
timestamp 1644511149
transform 1 0 30268 0 -1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_169_329
timestamp 1644511149
transform 1 0 31372 0 -1 94656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_169_335
timestamp 1644511149
transform 1 0 31924 0 -1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_169_337
timestamp 1644511149
transform 1 0 32108 0 -1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_169_349
timestamp 1644511149
transform 1 0 33212 0 -1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_169_361
timestamp 1644511149
transform 1 0 34316 0 -1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_169_373
timestamp 1644511149
transform 1 0 35420 0 -1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_169_385
timestamp 1644511149
transform 1 0 36524 0 -1 94656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_169_391
timestamp 1644511149
transform 1 0 37076 0 -1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_169_393
timestamp 1644511149
transform 1 0 37260 0 -1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_169_405
timestamp 1644511149
transform 1 0 38364 0 -1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_169_417
timestamp 1644511149
transform 1 0 39468 0 -1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_169_429
timestamp 1644511149
transform 1 0 40572 0 -1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_169_441
timestamp 1644511149
transform 1 0 41676 0 -1 94656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_169_447
timestamp 1644511149
transform 1 0 42228 0 -1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_169_449
timestamp 1644511149
transform 1 0 42412 0 -1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_169_461
timestamp 1644511149
transform 1 0 43516 0 -1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_169_473
timestamp 1644511149
transform 1 0 44620 0 -1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_169_485
timestamp 1644511149
transform 1 0 45724 0 -1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_169_497
timestamp 1644511149
transform 1 0 46828 0 -1 94656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_169_503
timestamp 1644511149
transform 1 0 47380 0 -1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_169_505
timestamp 1644511149
transform 1 0 47564 0 -1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_169_517
timestamp 1644511149
transform 1 0 48668 0 -1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_169_529
timestamp 1644511149
transform 1 0 49772 0 -1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_169_541
timestamp 1644511149
transform 1 0 50876 0 -1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_169_553
timestamp 1644511149
transform 1 0 51980 0 -1 94656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_169_559
timestamp 1644511149
transform 1 0 52532 0 -1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_169_561
timestamp 1644511149
transform 1 0 52716 0 -1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_169_573
timestamp 1644511149
transform 1 0 53820 0 -1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_169_585
timestamp 1644511149
transform 1 0 54924 0 -1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_169_597
timestamp 1644511149
transform 1 0 56028 0 -1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_169_609
timestamp 1644511149
transform 1 0 57132 0 -1 94656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_169_615
timestamp 1644511149
transform 1 0 57684 0 -1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_169_617
timestamp 1644511149
transform 1 0 57868 0 -1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_169_629
timestamp 1644511149
transform 1 0 58972 0 -1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_169_641
timestamp 1644511149
transform 1 0 60076 0 -1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_169_653
timestamp 1644511149
transform 1 0 61180 0 -1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_169_665
timestamp 1644511149
transform 1 0 62284 0 -1 94656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_169_671
timestamp 1644511149
transform 1 0 62836 0 -1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_169_673
timestamp 1644511149
transform 1 0 63020 0 -1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_169_685
timestamp 1644511149
transform 1 0 64124 0 -1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_169_697
timestamp 1644511149
transform 1 0 65228 0 -1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_169_709
timestamp 1644511149
transform 1 0 66332 0 -1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_169_721
timestamp 1644511149
transform 1 0 67436 0 -1 94656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_169_727
timestamp 1644511149
transform 1 0 67988 0 -1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_169_729
timestamp 1644511149
transform 1 0 68172 0 -1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_169_741
timestamp 1644511149
transform 1 0 69276 0 -1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_169_753
timestamp 1644511149
transform 1 0 70380 0 -1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_169_765
timestamp 1644511149
transform 1 0 71484 0 -1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_169_777
timestamp 1644511149
transform 1 0 72588 0 -1 94656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_169_783
timestamp 1644511149
transform 1 0 73140 0 -1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_169_785
timestamp 1644511149
transform 1 0 73324 0 -1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_169_797
timestamp 1644511149
transform 1 0 74428 0 -1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_169_809
timestamp 1644511149
transform 1 0 75532 0 -1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_169_821
timestamp 1644511149
transform 1 0 76636 0 -1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_169_833
timestamp 1644511149
transform 1 0 77740 0 -1 94656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_169_839
timestamp 1644511149
transform 1 0 78292 0 -1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_169_841
timestamp 1644511149
transform 1 0 78476 0 -1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_170_3
timestamp 1644511149
transform 1 0 1380 0 1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_170_15
timestamp 1644511149
transform 1 0 2484 0 1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_170_27
timestamp 1644511149
transform 1 0 3588 0 1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_170_29
timestamp 1644511149
transform 1 0 3772 0 1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_170_41
timestamp 1644511149
transform 1 0 4876 0 1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_170_53
timestamp 1644511149
transform 1 0 5980 0 1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_170_65
timestamp 1644511149
transform 1 0 7084 0 1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_170_77
timestamp 1644511149
transform 1 0 8188 0 1 94656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_170_83
timestamp 1644511149
transform 1 0 8740 0 1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_170_85
timestamp 1644511149
transform 1 0 8924 0 1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_170_97
timestamp 1644511149
transform 1 0 10028 0 1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_170_109
timestamp 1644511149
transform 1 0 11132 0 1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_170_121
timestamp 1644511149
transform 1 0 12236 0 1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_170_133
timestamp 1644511149
transform 1 0 13340 0 1 94656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_170_139
timestamp 1644511149
transform 1 0 13892 0 1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_170_141
timestamp 1644511149
transform 1 0 14076 0 1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_170_153
timestamp 1644511149
transform 1 0 15180 0 1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_170_165
timestamp 1644511149
transform 1 0 16284 0 1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_170_177
timestamp 1644511149
transform 1 0 17388 0 1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_170_189
timestamp 1644511149
transform 1 0 18492 0 1 94656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_170_195
timestamp 1644511149
transform 1 0 19044 0 1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_170_197
timestamp 1644511149
transform 1 0 19228 0 1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_170_209
timestamp 1644511149
transform 1 0 20332 0 1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_170_221
timestamp 1644511149
transform 1 0 21436 0 1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_170_233
timestamp 1644511149
transform 1 0 22540 0 1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_170_245
timestamp 1644511149
transform 1 0 23644 0 1 94656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_170_251
timestamp 1644511149
transform 1 0 24196 0 1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_170_253
timestamp 1644511149
transform 1 0 24380 0 1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_170_265
timestamp 1644511149
transform 1 0 25484 0 1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_170_277
timestamp 1644511149
transform 1 0 26588 0 1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_170_289
timestamp 1644511149
transform 1 0 27692 0 1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_170_301
timestamp 1644511149
transform 1 0 28796 0 1 94656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_170_307
timestamp 1644511149
transform 1 0 29348 0 1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_170_309
timestamp 1644511149
transform 1 0 29532 0 1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_170_321
timestamp 1644511149
transform 1 0 30636 0 1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_170_333
timestamp 1644511149
transform 1 0 31740 0 1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_170_345
timestamp 1644511149
transform 1 0 32844 0 1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_170_357
timestamp 1644511149
transform 1 0 33948 0 1 94656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_170_363
timestamp 1644511149
transform 1 0 34500 0 1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_170_365
timestamp 1644511149
transform 1 0 34684 0 1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_170_377
timestamp 1644511149
transform 1 0 35788 0 1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_170_389
timestamp 1644511149
transform 1 0 36892 0 1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_170_401
timestamp 1644511149
transform 1 0 37996 0 1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_170_413
timestamp 1644511149
transform 1 0 39100 0 1 94656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_170_419
timestamp 1644511149
transform 1 0 39652 0 1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_170_421
timestamp 1644511149
transform 1 0 39836 0 1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_170_433
timestamp 1644511149
transform 1 0 40940 0 1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_170_445
timestamp 1644511149
transform 1 0 42044 0 1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_170_457
timestamp 1644511149
transform 1 0 43148 0 1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_170_469
timestamp 1644511149
transform 1 0 44252 0 1 94656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_170_475
timestamp 1644511149
transform 1 0 44804 0 1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_170_477
timestamp 1644511149
transform 1 0 44988 0 1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_170_489
timestamp 1644511149
transform 1 0 46092 0 1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_170_501
timestamp 1644511149
transform 1 0 47196 0 1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_170_513
timestamp 1644511149
transform 1 0 48300 0 1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_170_525
timestamp 1644511149
transform 1 0 49404 0 1 94656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_170_531
timestamp 1644511149
transform 1 0 49956 0 1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_170_533
timestamp 1644511149
transform 1 0 50140 0 1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_170_545
timestamp 1644511149
transform 1 0 51244 0 1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_170_557
timestamp 1644511149
transform 1 0 52348 0 1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_170_569
timestamp 1644511149
transform 1 0 53452 0 1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_170_581
timestamp 1644511149
transform 1 0 54556 0 1 94656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_170_587
timestamp 1644511149
transform 1 0 55108 0 1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_170_589
timestamp 1644511149
transform 1 0 55292 0 1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_170_601
timestamp 1644511149
transform 1 0 56396 0 1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_170_613
timestamp 1644511149
transform 1 0 57500 0 1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_170_625
timestamp 1644511149
transform 1 0 58604 0 1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_170_637
timestamp 1644511149
transform 1 0 59708 0 1 94656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_170_643
timestamp 1644511149
transform 1 0 60260 0 1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_170_645
timestamp 1644511149
transform 1 0 60444 0 1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_170_657
timestamp 1644511149
transform 1 0 61548 0 1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_170_669
timestamp 1644511149
transform 1 0 62652 0 1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_170_681
timestamp 1644511149
transform 1 0 63756 0 1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_170_693
timestamp 1644511149
transform 1 0 64860 0 1 94656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_170_699
timestamp 1644511149
transform 1 0 65412 0 1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_170_701
timestamp 1644511149
transform 1 0 65596 0 1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_170_713
timestamp 1644511149
transform 1 0 66700 0 1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_170_725
timestamp 1644511149
transform 1 0 67804 0 1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_170_737
timestamp 1644511149
transform 1 0 68908 0 1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_170_749
timestamp 1644511149
transform 1 0 70012 0 1 94656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_170_755
timestamp 1644511149
transform 1 0 70564 0 1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_170_757
timestamp 1644511149
transform 1 0 70748 0 1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_170_769
timestamp 1644511149
transform 1 0 71852 0 1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_170_781
timestamp 1644511149
transform 1 0 72956 0 1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_170_793
timestamp 1644511149
transform 1 0 74060 0 1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_170_805
timestamp 1644511149
transform 1 0 75164 0 1 94656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_170_811
timestamp 1644511149
transform 1 0 75716 0 1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_170_813
timestamp 1644511149
transform 1 0 75900 0 1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_170_825
timestamp 1644511149
transform 1 0 77004 0 1 94656
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_170_833
timestamp 1644511149
transform 1 0 77740 0 1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_170_838
timestamp 1644511149
transform 1 0 78200 0 1 94656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_171_3
timestamp 1644511149
transform 1 0 1380 0 -1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_171_15
timestamp 1644511149
transform 1 0 2484 0 -1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_171_27
timestamp 1644511149
transform 1 0 3588 0 -1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_171_39
timestamp 1644511149
transform 1 0 4692 0 -1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_171_51
timestamp 1644511149
transform 1 0 5796 0 -1 95744
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_171_55
timestamp 1644511149
transform 1 0 6164 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_171_57
timestamp 1644511149
transform 1 0 6348 0 -1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_171_69
timestamp 1644511149
transform 1 0 7452 0 -1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_171_81
timestamp 1644511149
transform 1 0 8556 0 -1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_171_93
timestamp 1644511149
transform 1 0 9660 0 -1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_171_105
timestamp 1644511149
transform 1 0 10764 0 -1 95744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_171_111
timestamp 1644511149
transform 1 0 11316 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_171_113
timestamp 1644511149
transform 1 0 11500 0 -1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_171_125
timestamp 1644511149
transform 1 0 12604 0 -1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_171_137
timestamp 1644511149
transform 1 0 13708 0 -1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_171_149
timestamp 1644511149
transform 1 0 14812 0 -1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_171_161
timestamp 1644511149
transform 1 0 15916 0 -1 95744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_171_167
timestamp 1644511149
transform 1 0 16468 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_171_169
timestamp 1644511149
transform 1 0 16652 0 -1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_171_181
timestamp 1644511149
transform 1 0 17756 0 -1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_171_193
timestamp 1644511149
transform 1 0 18860 0 -1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_171_205
timestamp 1644511149
transform 1 0 19964 0 -1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_171_217
timestamp 1644511149
transform 1 0 21068 0 -1 95744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_171_223
timestamp 1644511149
transform 1 0 21620 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_171_225
timestamp 1644511149
transform 1 0 21804 0 -1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_171_237
timestamp 1644511149
transform 1 0 22908 0 -1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_171_249
timestamp 1644511149
transform 1 0 24012 0 -1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_171_261
timestamp 1644511149
transform 1 0 25116 0 -1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_171_273
timestamp 1644511149
transform 1 0 26220 0 -1 95744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_171_279
timestamp 1644511149
transform 1 0 26772 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_171_281
timestamp 1644511149
transform 1 0 26956 0 -1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_171_293
timestamp 1644511149
transform 1 0 28060 0 -1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_171_305
timestamp 1644511149
transform 1 0 29164 0 -1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_171_317
timestamp 1644511149
transform 1 0 30268 0 -1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_171_329
timestamp 1644511149
transform 1 0 31372 0 -1 95744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_171_335
timestamp 1644511149
transform 1 0 31924 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_171_337
timestamp 1644511149
transform 1 0 32108 0 -1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_171_349
timestamp 1644511149
transform 1 0 33212 0 -1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_171_361
timestamp 1644511149
transform 1 0 34316 0 -1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_171_373
timestamp 1644511149
transform 1 0 35420 0 -1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_171_385
timestamp 1644511149
transform 1 0 36524 0 -1 95744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_171_391
timestamp 1644511149
transform 1 0 37076 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_171_393
timestamp 1644511149
transform 1 0 37260 0 -1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_171_405
timestamp 1644511149
transform 1 0 38364 0 -1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_171_417
timestamp 1644511149
transform 1 0 39468 0 -1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_171_429
timestamp 1644511149
transform 1 0 40572 0 -1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_171_441
timestamp 1644511149
transform 1 0 41676 0 -1 95744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_171_447
timestamp 1644511149
transform 1 0 42228 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_171_449
timestamp 1644511149
transform 1 0 42412 0 -1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_171_461
timestamp 1644511149
transform 1 0 43516 0 -1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_171_473
timestamp 1644511149
transform 1 0 44620 0 -1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_171_485
timestamp 1644511149
transform 1 0 45724 0 -1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_171_497
timestamp 1644511149
transform 1 0 46828 0 -1 95744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_171_503
timestamp 1644511149
transform 1 0 47380 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_171_505
timestamp 1644511149
transform 1 0 47564 0 -1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_171_517
timestamp 1644511149
transform 1 0 48668 0 -1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_171_529
timestamp 1644511149
transform 1 0 49772 0 -1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_171_541
timestamp 1644511149
transform 1 0 50876 0 -1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_171_553
timestamp 1644511149
transform 1 0 51980 0 -1 95744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_171_559
timestamp 1644511149
transform 1 0 52532 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_171_561
timestamp 1644511149
transform 1 0 52716 0 -1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_171_573
timestamp 1644511149
transform 1 0 53820 0 -1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_171_585
timestamp 1644511149
transform 1 0 54924 0 -1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_171_597
timestamp 1644511149
transform 1 0 56028 0 -1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_171_609
timestamp 1644511149
transform 1 0 57132 0 -1 95744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_171_615
timestamp 1644511149
transform 1 0 57684 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_171_617
timestamp 1644511149
transform 1 0 57868 0 -1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_171_629
timestamp 1644511149
transform 1 0 58972 0 -1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_171_641
timestamp 1644511149
transform 1 0 60076 0 -1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_171_653
timestamp 1644511149
transform 1 0 61180 0 -1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_171_665
timestamp 1644511149
transform 1 0 62284 0 -1 95744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_171_671
timestamp 1644511149
transform 1 0 62836 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_171_673
timestamp 1644511149
transform 1 0 63020 0 -1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_171_685
timestamp 1644511149
transform 1 0 64124 0 -1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_171_697
timestamp 1644511149
transform 1 0 65228 0 -1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_171_709
timestamp 1644511149
transform 1 0 66332 0 -1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_171_721
timestamp 1644511149
transform 1 0 67436 0 -1 95744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_171_727
timestamp 1644511149
transform 1 0 67988 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_171_729
timestamp 1644511149
transform 1 0 68172 0 -1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_171_741
timestamp 1644511149
transform 1 0 69276 0 -1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_171_753
timestamp 1644511149
transform 1 0 70380 0 -1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_171_765
timestamp 1644511149
transform 1 0 71484 0 -1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_171_777
timestamp 1644511149
transform 1 0 72588 0 -1 95744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_171_783
timestamp 1644511149
transform 1 0 73140 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_171_785
timestamp 1644511149
transform 1 0 73324 0 -1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_171_797
timestamp 1644511149
transform 1 0 74428 0 -1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_171_809
timestamp 1644511149
transform 1 0 75532 0 -1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_171_821
timestamp 1644511149
transform 1 0 76636 0 -1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_171_833
timestamp 1644511149
transform 1 0 77740 0 -1 95744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_171_839
timestamp 1644511149
transform 1 0 78292 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_171_841
timestamp 1644511149
transform 1 0 78476 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_172_3
timestamp 1644511149
transform 1 0 1380 0 1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_172_15
timestamp 1644511149
transform 1 0 2484 0 1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_172_27
timestamp 1644511149
transform 1 0 3588 0 1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_172_29
timestamp 1644511149
transform 1 0 3772 0 1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_172_41
timestamp 1644511149
transform 1 0 4876 0 1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_172_53
timestamp 1644511149
transform 1 0 5980 0 1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_172_65
timestamp 1644511149
transform 1 0 7084 0 1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_172_77
timestamp 1644511149
transform 1 0 8188 0 1 95744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_172_83
timestamp 1644511149
transform 1 0 8740 0 1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_172_85
timestamp 1644511149
transform 1 0 8924 0 1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_172_97
timestamp 1644511149
transform 1 0 10028 0 1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_172_109
timestamp 1644511149
transform 1 0 11132 0 1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_172_121
timestamp 1644511149
transform 1 0 12236 0 1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_172_133
timestamp 1644511149
transform 1 0 13340 0 1 95744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_172_139
timestamp 1644511149
transform 1 0 13892 0 1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_172_141
timestamp 1644511149
transform 1 0 14076 0 1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_172_153
timestamp 1644511149
transform 1 0 15180 0 1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_172_165
timestamp 1644511149
transform 1 0 16284 0 1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_172_177
timestamp 1644511149
transform 1 0 17388 0 1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_172_189
timestamp 1644511149
transform 1 0 18492 0 1 95744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_172_195
timestamp 1644511149
transform 1 0 19044 0 1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_172_197
timestamp 1644511149
transform 1 0 19228 0 1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_172_209
timestamp 1644511149
transform 1 0 20332 0 1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_172_221
timestamp 1644511149
transform 1 0 21436 0 1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_172_233
timestamp 1644511149
transform 1 0 22540 0 1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_172_245
timestamp 1644511149
transform 1 0 23644 0 1 95744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_172_251
timestamp 1644511149
transform 1 0 24196 0 1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_172_253
timestamp 1644511149
transform 1 0 24380 0 1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_172_265
timestamp 1644511149
transform 1 0 25484 0 1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_172_277
timestamp 1644511149
transform 1 0 26588 0 1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_172_289
timestamp 1644511149
transform 1 0 27692 0 1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_172_301
timestamp 1644511149
transform 1 0 28796 0 1 95744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_172_307
timestamp 1644511149
transform 1 0 29348 0 1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_172_309
timestamp 1644511149
transform 1 0 29532 0 1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_172_321
timestamp 1644511149
transform 1 0 30636 0 1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_172_333
timestamp 1644511149
transform 1 0 31740 0 1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_172_345
timestamp 1644511149
transform 1 0 32844 0 1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_172_357
timestamp 1644511149
transform 1 0 33948 0 1 95744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_172_363
timestamp 1644511149
transform 1 0 34500 0 1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_172_365
timestamp 1644511149
transform 1 0 34684 0 1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_172_377
timestamp 1644511149
transform 1 0 35788 0 1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_172_389
timestamp 1644511149
transform 1 0 36892 0 1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_172_401
timestamp 1644511149
transform 1 0 37996 0 1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_172_413
timestamp 1644511149
transform 1 0 39100 0 1 95744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_172_419
timestamp 1644511149
transform 1 0 39652 0 1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_172_421
timestamp 1644511149
transform 1 0 39836 0 1 95744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_172_431
timestamp 1644511149
transform 1 0 40756 0 1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_172_443
timestamp 1644511149
transform 1 0 41860 0 1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_172_455
timestamp 1644511149
transform 1 0 42964 0 1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_172_467
timestamp 1644511149
transform 1 0 44068 0 1 95744
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_172_475
timestamp 1644511149
transform 1 0 44804 0 1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_172_477
timestamp 1644511149
transform 1 0 44988 0 1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_172_489
timestamp 1644511149
transform 1 0 46092 0 1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_172_501
timestamp 1644511149
transform 1 0 47196 0 1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_172_513
timestamp 1644511149
transform 1 0 48300 0 1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_172_525
timestamp 1644511149
transform 1 0 49404 0 1 95744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_172_531
timestamp 1644511149
transform 1 0 49956 0 1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_172_533
timestamp 1644511149
transform 1 0 50140 0 1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_172_545
timestamp 1644511149
transform 1 0 51244 0 1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_172_557
timestamp 1644511149
transform 1 0 52348 0 1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_172_569
timestamp 1644511149
transform 1 0 53452 0 1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_172_581
timestamp 1644511149
transform 1 0 54556 0 1 95744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_172_587
timestamp 1644511149
transform 1 0 55108 0 1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_172_589
timestamp 1644511149
transform 1 0 55292 0 1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_172_601
timestamp 1644511149
transform 1 0 56396 0 1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_172_613
timestamp 1644511149
transform 1 0 57500 0 1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_172_625
timestamp 1644511149
transform 1 0 58604 0 1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_172_637
timestamp 1644511149
transform 1 0 59708 0 1 95744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_172_643
timestamp 1644511149
transform 1 0 60260 0 1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_172_645
timestamp 1644511149
transform 1 0 60444 0 1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_172_657
timestamp 1644511149
transform 1 0 61548 0 1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_172_669
timestamp 1644511149
transform 1 0 62652 0 1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_172_681
timestamp 1644511149
transform 1 0 63756 0 1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_172_693
timestamp 1644511149
transform 1 0 64860 0 1 95744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_172_699
timestamp 1644511149
transform 1 0 65412 0 1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_172_701
timestamp 1644511149
transform 1 0 65596 0 1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_172_713
timestamp 1644511149
transform 1 0 66700 0 1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_172_725
timestamp 1644511149
transform 1 0 67804 0 1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_172_737
timestamp 1644511149
transform 1 0 68908 0 1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_172_749
timestamp 1644511149
transform 1 0 70012 0 1 95744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_172_755
timestamp 1644511149
transform 1 0 70564 0 1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_172_757
timestamp 1644511149
transform 1 0 70748 0 1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_172_769
timestamp 1644511149
transform 1 0 71852 0 1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_172_781
timestamp 1644511149
transform 1 0 72956 0 1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_172_793
timestamp 1644511149
transform 1 0 74060 0 1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_172_805
timestamp 1644511149
transform 1 0 75164 0 1 95744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_172_811
timestamp 1644511149
transform 1 0 75716 0 1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_172_813
timestamp 1644511149
transform 1 0 75900 0 1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_172_825
timestamp 1644511149
transform 1 0 77004 0 1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_172_837
timestamp 1644511149
transform 1 0 78108 0 1 95744
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_172_841
timestamp 1644511149
transform 1 0 78476 0 1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_173_3
timestamp 1644511149
transform 1 0 1380 0 -1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_173_15
timestamp 1644511149
transform 1 0 2484 0 -1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_173_27
timestamp 1644511149
transform 1 0 3588 0 -1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_173_39
timestamp 1644511149
transform 1 0 4692 0 -1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_173_51
timestamp 1644511149
transform 1 0 5796 0 -1 96832
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_173_55
timestamp 1644511149
transform 1 0 6164 0 -1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_173_57
timestamp 1644511149
transform 1 0 6348 0 -1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_173_69
timestamp 1644511149
transform 1 0 7452 0 -1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_173_81
timestamp 1644511149
transform 1 0 8556 0 -1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_173_93
timestamp 1644511149
transform 1 0 9660 0 -1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_173_105
timestamp 1644511149
transform 1 0 10764 0 -1 96832
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_173_111
timestamp 1644511149
transform 1 0 11316 0 -1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_173_113
timestamp 1644511149
transform 1 0 11500 0 -1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_173_125
timestamp 1644511149
transform 1 0 12604 0 -1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_173_137
timestamp 1644511149
transform 1 0 13708 0 -1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_173_149
timestamp 1644511149
transform 1 0 14812 0 -1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_173_161
timestamp 1644511149
transform 1 0 15916 0 -1 96832
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_173_167
timestamp 1644511149
transform 1 0 16468 0 -1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_173_169
timestamp 1644511149
transform 1 0 16652 0 -1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_173_181
timestamp 1644511149
transform 1 0 17756 0 -1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_173_193
timestamp 1644511149
transform 1 0 18860 0 -1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_173_205
timestamp 1644511149
transform 1 0 19964 0 -1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_173_217
timestamp 1644511149
transform 1 0 21068 0 -1 96832
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_173_223
timestamp 1644511149
transform 1 0 21620 0 -1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_173_225
timestamp 1644511149
transform 1 0 21804 0 -1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_173_237
timestamp 1644511149
transform 1 0 22908 0 -1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_173_249
timestamp 1644511149
transform 1 0 24012 0 -1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_173_261
timestamp 1644511149
transform 1 0 25116 0 -1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_173_273
timestamp 1644511149
transform 1 0 26220 0 -1 96832
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_173_279
timestamp 1644511149
transform 1 0 26772 0 -1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_173_281
timestamp 1644511149
transform 1 0 26956 0 -1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_173_293
timestamp 1644511149
transform 1 0 28060 0 -1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_173_305
timestamp 1644511149
transform 1 0 29164 0 -1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_173_317
timestamp 1644511149
transform 1 0 30268 0 -1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_173_329
timestamp 1644511149
transform 1 0 31372 0 -1 96832
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_173_335
timestamp 1644511149
transform 1 0 31924 0 -1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_173_337
timestamp 1644511149
transform 1 0 32108 0 -1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_173_349
timestamp 1644511149
transform 1 0 33212 0 -1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_173_361
timestamp 1644511149
transform 1 0 34316 0 -1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_173_373
timestamp 1644511149
transform 1 0 35420 0 -1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_173_385
timestamp 1644511149
transform 1 0 36524 0 -1 96832
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_173_391
timestamp 1644511149
transform 1 0 37076 0 -1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_173_393
timestamp 1644511149
transform 1 0 37260 0 -1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_173_405
timestamp 1644511149
transform 1 0 38364 0 -1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_173_417
timestamp 1644511149
transform 1 0 39468 0 -1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_173_429
timestamp 1644511149
transform 1 0 40572 0 -1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_173_441
timestamp 1644511149
transform 1 0 41676 0 -1 96832
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_173_447
timestamp 1644511149
transform 1 0 42228 0 -1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_173_449
timestamp 1644511149
transform 1 0 42412 0 -1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_173_461
timestamp 1644511149
transform 1 0 43516 0 -1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_173_473
timestamp 1644511149
transform 1 0 44620 0 -1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_173_485
timestamp 1644511149
transform 1 0 45724 0 -1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_173_497
timestamp 1644511149
transform 1 0 46828 0 -1 96832
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_173_503
timestamp 1644511149
transform 1 0 47380 0 -1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_173_505
timestamp 1644511149
transform 1 0 47564 0 -1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_173_517
timestamp 1644511149
transform 1 0 48668 0 -1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_173_529
timestamp 1644511149
transform 1 0 49772 0 -1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_173_541
timestamp 1644511149
transform 1 0 50876 0 -1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_173_553
timestamp 1644511149
transform 1 0 51980 0 -1 96832
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_173_559
timestamp 1644511149
transform 1 0 52532 0 -1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_173_561
timestamp 1644511149
transform 1 0 52716 0 -1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_173_573
timestamp 1644511149
transform 1 0 53820 0 -1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_173_585
timestamp 1644511149
transform 1 0 54924 0 -1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_173_597
timestamp 1644511149
transform 1 0 56028 0 -1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_173_609
timestamp 1644511149
transform 1 0 57132 0 -1 96832
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_173_615
timestamp 1644511149
transform 1 0 57684 0 -1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_173_617
timestamp 1644511149
transform 1 0 57868 0 -1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_173_629
timestamp 1644511149
transform 1 0 58972 0 -1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_173_641
timestamp 1644511149
transform 1 0 60076 0 -1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_173_653
timestamp 1644511149
transform 1 0 61180 0 -1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_173_665
timestamp 1644511149
transform 1 0 62284 0 -1 96832
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_173_671
timestamp 1644511149
transform 1 0 62836 0 -1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_173_673
timestamp 1644511149
transform 1 0 63020 0 -1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_173_685
timestamp 1644511149
transform 1 0 64124 0 -1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_173_697
timestamp 1644511149
transform 1 0 65228 0 -1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_173_709
timestamp 1644511149
transform 1 0 66332 0 -1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_173_721
timestamp 1644511149
transform 1 0 67436 0 -1 96832
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_173_727
timestamp 1644511149
transform 1 0 67988 0 -1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_173_729
timestamp 1644511149
transform 1 0 68172 0 -1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_173_741
timestamp 1644511149
transform 1 0 69276 0 -1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_173_753
timestamp 1644511149
transform 1 0 70380 0 -1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_173_765
timestamp 1644511149
transform 1 0 71484 0 -1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_173_777
timestamp 1644511149
transform 1 0 72588 0 -1 96832
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_173_783
timestamp 1644511149
transform 1 0 73140 0 -1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_173_785
timestamp 1644511149
transform 1 0 73324 0 -1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_173_797
timestamp 1644511149
transform 1 0 74428 0 -1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_173_809
timestamp 1644511149
transform 1 0 75532 0 -1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_173_821
timestamp 1644511149
transform 1 0 76636 0 -1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_173_833
timestamp 1644511149
transform 1 0 77740 0 -1 96832
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_173_839
timestamp 1644511149
transform 1 0 78292 0 -1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_173_841
timestamp 1644511149
transform 1 0 78476 0 -1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_174_3
timestamp 1644511149
transform 1 0 1380 0 1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_174_15
timestamp 1644511149
transform 1 0 2484 0 1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_174_27
timestamp 1644511149
transform 1 0 3588 0 1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_174_29
timestamp 1644511149
transform 1 0 3772 0 1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_174_41
timestamp 1644511149
transform 1 0 4876 0 1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_174_53
timestamp 1644511149
transform 1 0 5980 0 1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_174_65
timestamp 1644511149
transform 1 0 7084 0 1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_174_77
timestamp 1644511149
transform 1 0 8188 0 1 96832
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_174_83
timestamp 1644511149
transform 1 0 8740 0 1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_174_85
timestamp 1644511149
transform 1 0 8924 0 1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_174_97
timestamp 1644511149
transform 1 0 10028 0 1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_174_109
timestamp 1644511149
transform 1 0 11132 0 1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_174_121
timestamp 1644511149
transform 1 0 12236 0 1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_174_133
timestamp 1644511149
transform 1 0 13340 0 1 96832
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_174_139
timestamp 1644511149
transform 1 0 13892 0 1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_174_141
timestamp 1644511149
transform 1 0 14076 0 1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_174_153
timestamp 1644511149
transform 1 0 15180 0 1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_174_165
timestamp 1644511149
transform 1 0 16284 0 1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_174_177
timestamp 1644511149
transform 1 0 17388 0 1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_174_189
timestamp 1644511149
transform 1 0 18492 0 1 96832
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_174_195
timestamp 1644511149
transform 1 0 19044 0 1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_174_197
timestamp 1644511149
transform 1 0 19228 0 1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_174_209
timestamp 1644511149
transform 1 0 20332 0 1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_174_221
timestamp 1644511149
transform 1 0 21436 0 1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_174_233
timestamp 1644511149
transform 1 0 22540 0 1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_174_245
timestamp 1644511149
transform 1 0 23644 0 1 96832
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_174_251
timestamp 1644511149
transform 1 0 24196 0 1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_174_253
timestamp 1644511149
transform 1 0 24380 0 1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_174_265
timestamp 1644511149
transform 1 0 25484 0 1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_174_277
timestamp 1644511149
transform 1 0 26588 0 1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_174_289
timestamp 1644511149
transform 1 0 27692 0 1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_174_301
timestamp 1644511149
transform 1 0 28796 0 1 96832
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_174_307
timestamp 1644511149
transform 1 0 29348 0 1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_174_309
timestamp 1644511149
transform 1 0 29532 0 1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_174_321
timestamp 1644511149
transform 1 0 30636 0 1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_174_333
timestamp 1644511149
transform 1 0 31740 0 1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_174_345
timestamp 1644511149
transform 1 0 32844 0 1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_174_357
timestamp 1644511149
transform 1 0 33948 0 1 96832
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_174_363
timestamp 1644511149
transform 1 0 34500 0 1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_174_365
timestamp 1644511149
transform 1 0 34684 0 1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_174_377
timestamp 1644511149
transform 1 0 35788 0 1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_174_389
timestamp 1644511149
transform 1 0 36892 0 1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_174_401
timestamp 1644511149
transform 1 0 37996 0 1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_174_413
timestamp 1644511149
transform 1 0 39100 0 1 96832
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_174_419
timestamp 1644511149
transform 1 0 39652 0 1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_174_421
timestamp 1644511149
transform 1 0 39836 0 1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_174_433
timestamp 1644511149
transform 1 0 40940 0 1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_174_445
timestamp 1644511149
transform 1 0 42044 0 1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_174_457
timestamp 1644511149
transform 1 0 43148 0 1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_174_469
timestamp 1644511149
transform 1 0 44252 0 1 96832
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_174_475
timestamp 1644511149
transform 1 0 44804 0 1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_174_477
timestamp 1644511149
transform 1 0 44988 0 1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_174_489
timestamp 1644511149
transform 1 0 46092 0 1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_174_501
timestamp 1644511149
transform 1 0 47196 0 1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_174_513
timestamp 1644511149
transform 1 0 48300 0 1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_174_525
timestamp 1644511149
transform 1 0 49404 0 1 96832
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_174_531
timestamp 1644511149
transform 1 0 49956 0 1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_174_533
timestamp 1644511149
transform 1 0 50140 0 1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_174_545
timestamp 1644511149
transform 1 0 51244 0 1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_174_557
timestamp 1644511149
transform 1 0 52348 0 1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_174_569
timestamp 1644511149
transform 1 0 53452 0 1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_174_581
timestamp 1644511149
transform 1 0 54556 0 1 96832
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_174_587
timestamp 1644511149
transform 1 0 55108 0 1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_174_589
timestamp 1644511149
transform 1 0 55292 0 1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_174_601
timestamp 1644511149
transform 1 0 56396 0 1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_174_613
timestamp 1644511149
transform 1 0 57500 0 1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_174_625
timestamp 1644511149
transform 1 0 58604 0 1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_174_637
timestamp 1644511149
transform 1 0 59708 0 1 96832
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_174_643
timestamp 1644511149
transform 1 0 60260 0 1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_174_645
timestamp 1644511149
transform 1 0 60444 0 1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_174_657
timestamp 1644511149
transform 1 0 61548 0 1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_174_669
timestamp 1644511149
transform 1 0 62652 0 1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_174_681
timestamp 1644511149
transform 1 0 63756 0 1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_174_693
timestamp 1644511149
transform 1 0 64860 0 1 96832
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_174_699
timestamp 1644511149
transform 1 0 65412 0 1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_174_701
timestamp 1644511149
transform 1 0 65596 0 1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_174_713
timestamp 1644511149
transform 1 0 66700 0 1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_174_725
timestamp 1644511149
transform 1 0 67804 0 1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_174_737
timestamp 1644511149
transform 1 0 68908 0 1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_174_749
timestamp 1644511149
transform 1 0 70012 0 1 96832
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_174_755
timestamp 1644511149
transform 1 0 70564 0 1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_174_757
timestamp 1644511149
transform 1 0 70748 0 1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_174_769
timestamp 1644511149
transform 1 0 71852 0 1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_174_781
timestamp 1644511149
transform 1 0 72956 0 1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_174_793
timestamp 1644511149
transform 1 0 74060 0 1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_174_805
timestamp 1644511149
transform 1 0 75164 0 1 96832
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_174_811
timestamp 1644511149
transform 1 0 75716 0 1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_174_813
timestamp 1644511149
transform 1 0 75900 0 1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_174_825
timestamp 1644511149
transform 1 0 77004 0 1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_174_837
timestamp 1644511149
transform 1 0 78108 0 1 96832
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_174_841
timestamp 1644511149
transform 1 0 78476 0 1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_175_9
timestamp 1644511149
transform 1 0 1932 0 -1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_175_21
timestamp 1644511149
transform 1 0 3036 0 -1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_175_33
timestamp 1644511149
transform 1 0 4140 0 -1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_175_45
timestamp 1644511149
transform 1 0 5244 0 -1 97920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_175_53
timestamp 1644511149
transform 1 0 5980 0 -1 97920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_175_57
timestamp 1644511149
transform 1 0 6348 0 -1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_175_69
timestamp 1644511149
transform 1 0 7452 0 -1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_175_81
timestamp 1644511149
transform 1 0 8556 0 -1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_175_93
timestamp 1644511149
transform 1 0 9660 0 -1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_175_105
timestamp 1644511149
transform 1 0 10764 0 -1 97920
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_175_111
timestamp 1644511149
transform 1 0 11316 0 -1 97920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_175_113
timestamp 1644511149
transform 1 0 11500 0 -1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_175_125
timestamp 1644511149
transform 1 0 12604 0 -1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_175_137
timestamp 1644511149
transform 1 0 13708 0 -1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_175_149
timestamp 1644511149
transform 1 0 14812 0 -1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_175_161
timestamp 1644511149
transform 1 0 15916 0 -1 97920
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_175_167
timestamp 1644511149
transform 1 0 16468 0 -1 97920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_175_169
timestamp 1644511149
transform 1 0 16652 0 -1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_175_181
timestamp 1644511149
transform 1 0 17756 0 -1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_175_193
timestamp 1644511149
transform 1 0 18860 0 -1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_175_205
timestamp 1644511149
transform 1 0 19964 0 -1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_175_217
timestamp 1644511149
transform 1 0 21068 0 -1 97920
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_175_223
timestamp 1644511149
transform 1 0 21620 0 -1 97920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_175_225
timestamp 1644511149
transform 1 0 21804 0 -1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_175_237
timestamp 1644511149
transform 1 0 22908 0 -1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_175_249
timestamp 1644511149
transform 1 0 24012 0 -1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_175_261
timestamp 1644511149
transform 1 0 25116 0 -1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_175_273
timestamp 1644511149
transform 1 0 26220 0 -1 97920
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_175_279
timestamp 1644511149
transform 1 0 26772 0 -1 97920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_175_281
timestamp 1644511149
transform 1 0 26956 0 -1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_175_293
timestamp 1644511149
transform 1 0 28060 0 -1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_175_305
timestamp 1644511149
transform 1 0 29164 0 -1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_175_317
timestamp 1644511149
transform 1 0 30268 0 -1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_175_329
timestamp 1644511149
transform 1 0 31372 0 -1 97920
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_175_335
timestamp 1644511149
transform 1 0 31924 0 -1 97920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_175_337
timestamp 1644511149
transform 1 0 32108 0 -1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_175_349
timestamp 1644511149
transform 1 0 33212 0 -1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_175_361
timestamp 1644511149
transform 1 0 34316 0 -1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_175_373
timestamp 1644511149
transform 1 0 35420 0 -1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_175_385
timestamp 1644511149
transform 1 0 36524 0 -1 97920
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_175_391
timestamp 1644511149
transform 1 0 37076 0 -1 97920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_175_393
timestamp 1644511149
transform 1 0 37260 0 -1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_175_405
timestamp 1644511149
transform 1 0 38364 0 -1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_175_417
timestamp 1644511149
transform 1 0 39468 0 -1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_175_429
timestamp 1644511149
transform 1 0 40572 0 -1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_175_441
timestamp 1644511149
transform 1 0 41676 0 -1 97920
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_175_447
timestamp 1644511149
transform 1 0 42228 0 -1 97920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_175_449
timestamp 1644511149
transform 1 0 42412 0 -1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_175_461
timestamp 1644511149
transform 1 0 43516 0 -1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_175_473
timestamp 1644511149
transform 1 0 44620 0 -1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_175_485
timestamp 1644511149
transform 1 0 45724 0 -1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_175_497
timestamp 1644511149
transform 1 0 46828 0 -1 97920
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_175_503
timestamp 1644511149
transform 1 0 47380 0 -1 97920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_175_505
timestamp 1644511149
transform 1 0 47564 0 -1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_175_517
timestamp 1644511149
transform 1 0 48668 0 -1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_175_529
timestamp 1644511149
transform 1 0 49772 0 -1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_175_541
timestamp 1644511149
transform 1 0 50876 0 -1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_175_553
timestamp 1644511149
transform 1 0 51980 0 -1 97920
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_175_559
timestamp 1644511149
transform 1 0 52532 0 -1 97920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_175_561
timestamp 1644511149
transform 1 0 52716 0 -1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_175_573
timestamp 1644511149
transform 1 0 53820 0 -1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_175_585
timestamp 1644511149
transform 1 0 54924 0 -1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_175_597
timestamp 1644511149
transform 1 0 56028 0 -1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_175_609
timestamp 1644511149
transform 1 0 57132 0 -1 97920
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_175_615
timestamp 1644511149
transform 1 0 57684 0 -1 97920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_175_617
timestamp 1644511149
transform 1 0 57868 0 -1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_175_629
timestamp 1644511149
transform 1 0 58972 0 -1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_175_641
timestamp 1644511149
transform 1 0 60076 0 -1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_175_653
timestamp 1644511149
transform 1 0 61180 0 -1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_175_665
timestamp 1644511149
transform 1 0 62284 0 -1 97920
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_175_671
timestamp 1644511149
transform 1 0 62836 0 -1 97920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_175_673
timestamp 1644511149
transform 1 0 63020 0 -1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_175_685
timestamp 1644511149
transform 1 0 64124 0 -1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_175_697
timestamp 1644511149
transform 1 0 65228 0 -1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_175_709
timestamp 1644511149
transform 1 0 66332 0 -1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_175_721
timestamp 1644511149
transform 1 0 67436 0 -1 97920
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_175_727
timestamp 1644511149
transform 1 0 67988 0 -1 97920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_175_729
timestamp 1644511149
transform 1 0 68172 0 -1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_175_741
timestamp 1644511149
transform 1 0 69276 0 -1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_175_753
timestamp 1644511149
transform 1 0 70380 0 -1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_175_765
timestamp 1644511149
transform 1 0 71484 0 -1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_175_777
timestamp 1644511149
transform 1 0 72588 0 -1 97920
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_175_783
timestamp 1644511149
transform 1 0 73140 0 -1 97920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_175_785
timestamp 1644511149
transform 1 0 73324 0 -1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_175_797
timestamp 1644511149
transform 1 0 74428 0 -1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_175_809
timestamp 1644511149
transform 1 0 75532 0 -1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_175_821
timestamp 1644511149
transform 1 0 76636 0 -1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_175_833
timestamp 1644511149
transform 1 0 77740 0 -1 97920
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_175_839
timestamp 1644511149
transform 1 0 78292 0 -1 97920
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_175_841
timestamp 1644511149
transform 1 0 78476 0 -1 97920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_176_3
timestamp 1644511149
transform 1 0 1380 0 1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_176_15
timestamp 1644511149
transform 1 0 2484 0 1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_176_27
timestamp 1644511149
transform 1 0 3588 0 1 97920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_176_29
timestamp 1644511149
transform 1 0 3772 0 1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_176_41
timestamp 1644511149
transform 1 0 4876 0 1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_176_53
timestamp 1644511149
transform 1 0 5980 0 1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_176_65
timestamp 1644511149
transform 1 0 7084 0 1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_176_77
timestamp 1644511149
transform 1 0 8188 0 1 97920
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_176_83
timestamp 1644511149
transform 1 0 8740 0 1 97920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_176_85
timestamp 1644511149
transform 1 0 8924 0 1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_176_97
timestamp 1644511149
transform 1 0 10028 0 1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_176_109
timestamp 1644511149
transform 1 0 11132 0 1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_176_121
timestamp 1644511149
transform 1 0 12236 0 1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_176_133
timestamp 1644511149
transform 1 0 13340 0 1 97920
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_176_139
timestamp 1644511149
transform 1 0 13892 0 1 97920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_176_141
timestamp 1644511149
transform 1 0 14076 0 1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_176_153
timestamp 1644511149
transform 1 0 15180 0 1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_176_165
timestamp 1644511149
transform 1 0 16284 0 1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_176_177
timestamp 1644511149
transform 1 0 17388 0 1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_176_189
timestamp 1644511149
transform 1 0 18492 0 1 97920
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_176_195
timestamp 1644511149
transform 1 0 19044 0 1 97920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_176_197
timestamp 1644511149
transform 1 0 19228 0 1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_176_209
timestamp 1644511149
transform 1 0 20332 0 1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_176_221
timestamp 1644511149
transform 1 0 21436 0 1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_176_233
timestamp 1644511149
transform 1 0 22540 0 1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_176_245
timestamp 1644511149
transform 1 0 23644 0 1 97920
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_176_251
timestamp 1644511149
transform 1 0 24196 0 1 97920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_176_253
timestamp 1644511149
transform 1 0 24380 0 1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_176_265
timestamp 1644511149
transform 1 0 25484 0 1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_176_277
timestamp 1644511149
transform 1 0 26588 0 1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_176_289
timestamp 1644511149
transform 1 0 27692 0 1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_176_301
timestamp 1644511149
transform 1 0 28796 0 1 97920
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_176_307
timestamp 1644511149
transform 1 0 29348 0 1 97920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_176_309
timestamp 1644511149
transform 1 0 29532 0 1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_176_321
timestamp 1644511149
transform 1 0 30636 0 1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_176_333
timestamp 1644511149
transform 1 0 31740 0 1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_176_345
timestamp 1644511149
transform 1 0 32844 0 1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_176_357
timestamp 1644511149
transform 1 0 33948 0 1 97920
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_176_363
timestamp 1644511149
transform 1 0 34500 0 1 97920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_176_365
timestamp 1644511149
transform 1 0 34684 0 1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_176_377
timestamp 1644511149
transform 1 0 35788 0 1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_176_389
timestamp 1644511149
transform 1 0 36892 0 1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_176_401
timestamp 1644511149
transform 1 0 37996 0 1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_176_413
timestamp 1644511149
transform 1 0 39100 0 1 97920
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_176_419
timestamp 1644511149
transform 1 0 39652 0 1 97920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_176_421
timestamp 1644511149
transform 1 0 39836 0 1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_176_433
timestamp 1644511149
transform 1 0 40940 0 1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_176_445
timestamp 1644511149
transform 1 0 42044 0 1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_176_457
timestamp 1644511149
transform 1 0 43148 0 1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_176_469
timestamp 1644511149
transform 1 0 44252 0 1 97920
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_176_475
timestamp 1644511149
transform 1 0 44804 0 1 97920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_176_477
timestamp 1644511149
transform 1 0 44988 0 1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_176_489
timestamp 1644511149
transform 1 0 46092 0 1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_176_501
timestamp 1644511149
transform 1 0 47196 0 1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_176_513
timestamp 1644511149
transform 1 0 48300 0 1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_176_525
timestamp 1644511149
transform 1 0 49404 0 1 97920
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_176_531
timestamp 1644511149
transform 1 0 49956 0 1 97920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_176_533
timestamp 1644511149
transform 1 0 50140 0 1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_176_545
timestamp 1644511149
transform 1 0 51244 0 1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_176_557
timestamp 1644511149
transform 1 0 52348 0 1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_176_569
timestamp 1644511149
transform 1 0 53452 0 1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_176_581
timestamp 1644511149
transform 1 0 54556 0 1 97920
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_176_587
timestamp 1644511149
transform 1 0 55108 0 1 97920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_176_589
timestamp 1644511149
transform 1 0 55292 0 1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_176_601
timestamp 1644511149
transform 1 0 56396 0 1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_176_613
timestamp 1644511149
transform 1 0 57500 0 1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_176_625
timestamp 1644511149
transform 1 0 58604 0 1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_176_637
timestamp 1644511149
transform 1 0 59708 0 1 97920
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_176_643
timestamp 1644511149
transform 1 0 60260 0 1 97920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_176_645
timestamp 1644511149
transform 1 0 60444 0 1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_176_657
timestamp 1644511149
transform 1 0 61548 0 1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_176_669
timestamp 1644511149
transform 1 0 62652 0 1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_176_681
timestamp 1644511149
transform 1 0 63756 0 1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_176_693
timestamp 1644511149
transform 1 0 64860 0 1 97920
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_176_699
timestamp 1644511149
transform 1 0 65412 0 1 97920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_176_701
timestamp 1644511149
transform 1 0 65596 0 1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_176_713
timestamp 1644511149
transform 1 0 66700 0 1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_176_725
timestamp 1644511149
transform 1 0 67804 0 1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_176_737
timestamp 1644511149
transform 1 0 68908 0 1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_176_749
timestamp 1644511149
transform 1 0 70012 0 1 97920
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_176_755
timestamp 1644511149
transform 1 0 70564 0 1 97920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_176_757
timestamp 1644511149
transform 1 0 70748 0 1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_176_769
timestamp 1644511149
transform 1 0 71852 0 1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_176_781
timestamp 1644511149
transform 1 0 72956 0 1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_176_793
timestamp 1644511149
transform 1 0 74060 0 1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_176_805
timestamp 1644511149
transform 1 0 75164 0 1 97920
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_176_811
timestamp 1644511149
transform 1 0 75716 0 1 97920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_176_813
timestamp 1644511149
transform 1 0 75900 0 1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_176_825
timestamp 1644511149
transform 1 0 77004 0 1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_176_837
timestamp 1644511149
transform 1 0 78108 0 1 97920
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_176_841
timestamp 1644511149
transform 1 0 78476 0 1 97920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_177_3
timestamp 1644511149
transform 1 0 1380 0 -1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_177_15
timestamp 1644511149
transform 1 0 2484 0 -1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_177_27
timestamp 1644511149
transform 1 0 3588 0 -1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_177_39
timestamp 1644511149
transform 1 0 4692 0 -1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_177_51
timestamp 1644511149
transform 1 0 5796 0 -1 99008
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_177_55
timestamp 1644511149
transform 1 0 6164 0 -1 99008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_177_57
timestamp 1644511149
transform 1 0 6348 0 -1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_177_69
timestamp 1644511149
transform 1 0 7452 0 -1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_177_81
timestamp 1644511149
transform 1 0 8556 0 -1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_177_93
timestamp 1644511149
transform 1 0 9660 0 -1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_177_105
timestamp 1644511149
transform 1 0 10764 0 -1 99008
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_177_111
timestamp 1644511149
transform 1 0 11316 0 -1 99008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_177_113
timestamp 1644511149
transform 1 0 11500 0 -1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_177_125
timestamp 1644511149
transform 1 0 12604 0 -1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_177_137
timestamp 1644511149
transform 1 0 13708 0 -1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_177_149
timestamp 1644511149
transform 1 0 14812 0 -1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_177_161
timestamp 1644511149
transform 1 0 15916 0 -1 99008
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_177_167
timestamp 1644511149
transform 1 0 16468 0 -1 99008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_177_169
timestamp 1644511149
transform 1 0 16652 0 -1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_177_181
timestamp 1644511149
transform 1 0 17756 0 -1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_177_193
timestamp 1644511149
transform 1 0 18860 0 -1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_177_205
timestamp 1644511149
transform 1 0 19964 0 -1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_177_217
timestamp 1644511149
transform 1 0 21068 0 -1 99008
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_177_223
timestamp 1644511149
transform 1 0 21620 0 -1 99008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_177_225
timestamp 1644511149
transform 1 0 21804 0 -1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_177_237
timestamp 1644511149
transform 1 0 22908 0 -1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_177_249
timestamp 1644511149
transform 1 0 24012 0 -1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_177_261
timestamp 1644511149
transform 1 0 25116 0 -1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_177_273
timestamp 1644511149
transform 1 0 26220 0 -1 99008
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_177_279
timestamp 1644511149
transform 1 0 26772 0 -1 99008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_177_281
timestamp 1644511149
transform 1 0 26956 0 -1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_177_293
timestamp 1644511149
transform 1 0 28060 0 -1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_177_305
timestamp 1644511149
transform 1 0 29164 0 -1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_177_317
timestamp 1644511149
transform 1 0 30268 0 -1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_177_329
timestamp 1644511149
transform 1 0 31372 0 -1 99008
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_177_335
timestamp 1644511149
transform 1 0 31924 0 -1 99008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_177_337
timestamp 1644511149
transform 1 0 32108 0 -1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_177_349
timestamp 1644511149
transform 1 0 33212 0 -1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_177_361
timestamp 1644511149
transform 1 0 34316 0 -1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_177_373
timestamp 1644511149
transform 1 0 35420 0 -1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_177_385
timestamp 1644511149
transform 1 0 36524 0 -1 99008
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_177_391
timestamp 1644511149
transform 1 0 37076 0 -1 99008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_177_393
timestamp 1644511149
transform 1 0 37260 0 -1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_177_405
timestamp 1644511149
transform 1 0 38364 0 -1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_177_417
timestamp 1644511149
transform 1 0 39468 0 -1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_177_429
timestamp 1644511149
transform 1 0 40572 0 -1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_177_441
timestamp 1644511149
transform 1 0 41676 0 -1 99008
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_177_447
timestamp 1644511149
transform 1 0 42228 0 -1 99008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_177_449
timestamp 1644511149
transform 1 0 42412 0 -1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_177_461
timestamp 1644511149
transform 1 0 43516 0 -1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_177_473
timestamp 1644511149
transform 1 0 44620 0 -1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_177_485
timestamp 1644511149
transform 1 0 45724 0 -1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_177_497
timestamp 1644511149
transform 1 0 46828 0 -1 99008
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_177_503
timestamp 1644511149
transform 1 0 47380 0 -1 99008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_177_505
timestamp 1644511149
transform 1 0 47564 0 -1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_177_517
timestamp 1644511149
transform 1 0 48668 0 -1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_177_529
timestamp 1644511149
transform 1 0 49772 0 -1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_177_541
timestamp 1644511149
transform 1 0 50876 0 -1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_177_553
timestamp 1644511149
transform 1 0 51980 0 -1 99008
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_177_559
timestamp 1644511149
transform 1 0 52532 0 -1 99008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_177_561
timestamp 1644511149
transform 1 0 52716 0 -1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_177_573
timestamp 1644511149
transform 1 0 53820 0 -1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_177_585
timestamp 1644511149
transform 1 0 54924 0 -1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_177_597
timestamp 1644511149
transform 1 0 56028 0 -1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_177_609
timestamp 1644511149
transform 1 0 57132 0 -1 99008
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_177_615
timestamp 1644511149
transform 1 0 57684 0 -1 99008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_177_617
timestamp 1644511149
transform 1 0 57868 0 -1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_177_629
timestamp 1644511149
transform 1 0 58972 0 -1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_177_641
timestamp 1644511149
transform 1 0 60076 0 -1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_177_653
timestamp 1644511149
transform 1 0 61180 0 -1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_177_665
timestamp 1644511149
transform 1 0 62284 0 -1 99008
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_177_671
timestamp 1644511149
transform 1 0 62836 0 -1 99008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_177_673
timestamp 1644511149
transform 1 0 63020 0 -1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_177_685
timestamp 1644511149
transform 1 0 64124 0 -1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_177_697
timestamp 1644511149
transform 1 0 65228 0 -1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_177_709
timestamp 1644511149
transform 1 0 66332 0 -1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_177_721
timestamp 1644511149
transform 1 0 67436 0 -1 99008
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_177_727
timestamp 1644511149
transform 1 0 67988 0 -1 99008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_177_729
timestamp 1644511149
transform 1 0 68172 0 -1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_177_741
timestamp 1644511149
transform 1 0 69276 0 -1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_177_753
timestamp 1644511149
transform 1 0 70380 0 -1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_177_765
timestamp 1644511149
transform 1 0 71484 0 -1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_177_777
timestamp 1644511149
transform 1 0 72588 0 -1 99008
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_177_783
timestamp 1644511149
transform 1 0 73140 0 -1 99008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_177_785
timestamp 1644511149
transform 1 0 73324 0 -1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_177_797
timestamp 1644511149
transform 1 0 74428 0 -1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_177_809
timestamp 1644511149
transform 1 0 75532 0 -1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_177_821
timestamp 1644511149
transform 1 0 76636 0 -1 99008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_177_829
timestamp 1644511149
transform 1 0 77372 0 -1 99008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_177_836
timestamp 1644511149
transform 1 0 78016 0 -1 99008
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_177_841
timestamp 1644511149
transform 1 0 78476 0 -1 99008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_178_3
timestamp 1644511149
transform 1 0 1380 0 1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_178_15
timestamp 1644511149
transform 1 0 2484 0 1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_178_27
timestamp 1644511149
transform 1 0 3588 0 1 99008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_178_29
timestamp 1644511149
transform 1 0 3772 0 1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_178_41
timestamp 1644511149
transform 1 0 4876 0 1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_178_53
timestamp 1644511149
transform 1 0 5980 0 1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_178_65
timestamp 1644511149
transform 1 0 7084 0 1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_178_77
timestamp 1644511149
transform 1 0 8188 0 1 99008
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_178_83
timestamp 1644511149
transform 1 0 8740 0 1 99008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_178_85
timestamp 1644511149
transform 1 0 8924 0 1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_178_97
timestamp 1644511149
transform 1 0 10028 0 1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_178_109
timestamp 1644511149
transform 1 0 11132 0 1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_178_121
timestamp 1644511149
transform 1 0 12236 0 1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_178_133
timestamp 1644511149
transform 1 0 13340 0 1 99008
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_178_139
timestamp 1644511149
transform 1 0 13892 0 1 99008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_178_141
timestamp 1644511149
transform 1 0 14076 0 1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_178_153
timestamp 1644511149
transform 1 0 15180 0 1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_178_165
timestamp 1644511149
transform 1 0 16284 0 1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_178_177
timestamp 1644511149
transform 1 0 17388 0 1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_178_189
timestamp 1644511149
transform 1 0 18492 0 1 99008
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_178_195
timestamp 1644511149
transform 1 0 19044 0 1 99008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_178_197
timestamp 1644511149
transform 1 0 19228 0 1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_178_209
timestamp 1644511149
transform 1 0 20332 0 1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_178_221
timestamp 1644511149
transform 1 0 21436 0 1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_178_233
timestamp 1644511149
transform 1 0 22540 0 1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_178_245
timestamp 1644511149
transform 1 0 23644 0 1 99008
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_178_251
timestamp 1644511149
transform 1 0 24196 0 1 99008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_178_253
timestamp 1644511149
transform 1 0 24380 0 1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_178_265
timestamp 1644511149
transform 1 0 25484 0 1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_178_277
timestamp 1644511149
transform 1 0 26588 0 1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_178_289
timestamp 1644511149
transform 1 0 27692 0 1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_178_301
timestamp 1644511149
transform 1 0 28796 0 1 99008
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_178_307
timestamp 1644511149
transform 1 0 29348 0 1 99008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_178_309
timestamp 1644511149
transform 1 0 29532 0 1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_178_321
timestamp 1644511149
transform 1 0 30636 0 1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_178_333
timestamp 1644511149
transform 1 0 31740 0 1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_178_345
timestamp 1644511149
transform 1 0 32844 0 1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_178_357
timestamp 1644511149
transform 1 0 33948 0 1 99008
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_178_363
timestamp 1644511149
transform 1 0 34500 0 1 99008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_178_365
timestamp 1644511149
transform 1 0 34684 0 1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_178_377
timestamp 1644511149
transform 1 0 35788 0 1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_178_389
timestamp 1644511149
transform 1 0 36892 0 1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_178_401
timestamp 1644511149
transform 1 0 37996 0 1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_178_413
timestamp 1644511149
transform 1 0 39100 0 1 99008
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_178_419
timestamp 1644511149
transform 1 0 39652 0 1 99008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_178_421
timestamp 1644511149
transform 1 0 39836 0 1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_178_433
timestamp 1644511149
transform 1 0 40940 0 1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_178_445
timestamp 1644511149
transform 1 0 42044 0 1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_178_457
timestamp 1644511149
transform 1 0 43148 0 1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_178_469
timestamp 1644511149
transform 1 0 44252 0 1 99008
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_178_475
timestamp 1644511149
transform 1 0 44804 0 1 99008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_178_477
timestamp 1644511149
transform 1 0 44988 0 1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_178_489
timestamp 1644511149
transform 1 0 46092 0 1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_178_501
timestamp 1644511149
transform 1 0 47196 0 1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_178_513
timestamp 1644511149
transform 1 0 48300 0 1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_178_525
timestamp 1644511149
transform 1 0 49404 0 1 99008
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_178_531
timestamp 1644511149
transform 1 0 49956 0 1 99008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_178_533
timestamp 1644511149
transform 1 0 50140 0 1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_178_545
timestamp 1644511149
transform 1 0 51244 0 1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_178_557
timestamp 1644511149
transform 1 0 52348 0 1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_178_569
timestamp 1644511149
transform 1 0 53452 0 1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_178_581
timestamp 1644511149
transform 1 0 54556 0 1 99008
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_178_587
timestamp 1644511149
transform 1 0 55108 0 1 99008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_178_589
timestamp 1644511149
transform 1 0 55292 0 1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_178_601
timestamp 1644511149
transform 1 0 56396 0 1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_178_613
timestamp 1644511149
transform 1 0 57500 0 1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_178_625
timestamp 1644511149
transform 1 0 58604 0 1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_178_637
timestamp 1644511149
transform 1 0 59708 0 1 99008
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_178_643
timestamp 1644511149
transform 1 0 60260 0 1 99008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_178_645
timestamp 1644511149
transform 1 0 60444 0 1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_178_657
timestamp 1644511149
transform 1 0 61548 0 1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_178_669
timestamp 1644511149
transform 1 0 62652 0 1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_178_681
timestamp 1644511149
transform 1 0 63756 0 1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_178_693
timestamp 1644511149
transform 1 0 64860 0 1 99008
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_178_699
timestamp 1644511149
transform 1 0 65412 0 1 99008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_178_701
timestamp 1644511149
transform 1 0 65596 0 1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_178_713
timestamp 1644511149
transform 1 0 66700 0 1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_178_725
timestamp 1644511149
transform 1 0 67804 0 1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_178_737
timestamp 1644511149
transform 1 0 68908 0 1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_178_749
timestamp 1644511149
transform 1 0 70012 0 1 99008
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_178_755
timestamp 1644511149
transform 1 0 70564 0 1 99008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_178_757
timestamp 1644511149
transform 1 0 70748 0 1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_178_769
timestamp 1644511149
transform 1 0 71852 0 1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_178_781
timestamp 1644511149
transform 1 0 72956 0 1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_178_793
timestamp 1644511149
transform 1 0 74060 0 1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_178_805
timestamp 1644511149
transform 1 0 75164 0 1 99008
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_178_811
timestamp 1644511149
transform 1 0 75716 0 1 99008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_178_813
timestamp 1644511149
transform 1 0 75900 0 1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_178_825
timestamp 1644511149
transform 1 0 77004 0 1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_178_837
timestamp 1644511149
transform 1 0 78108 0 1 99008
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_178_841
timestamp 1644511149
transform 1 0 78476 0 1 99008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_179_3
timestamp 1644511149
transform 1 0 1380 0 -1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_179_15
timestamp 1644511149
transform 1 0 2484 0 -1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_179_27
timestamp 1644511149
transform 1 0 3588 0 -1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_179_39
timestamp 1644511149
transform 1 0 4692 0 -1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_179_51
timestamp 1644511149
transform 1 0 5796 0 -1 100096
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_179_55
timestamp 1644511149
transform 1 0 6164 0 -1 100096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_179_57
timestamp 1644511149
transform 1 0 6348 0 -1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_179_69
timestamp 1644511149
transform 1 0 7452 0 -1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_179_81
timestamp 1644511149
transform 1 0 8556 0 -1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_179_93
timestamp 1644511149
transform 1 0 9660 0 -1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_179_105
timestamp 1644511149
transform 1 0 10764 0 -1 100096
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_179_111
timestamp 1644511149
transform 1 0 11316 0 -1 100096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_179_113
timestamp 1644511149
transform 1 0 11500 0 -1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_179_125
timestamp 1644511149
transform 1 0 12604 0 -1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_179_137
timestamp 1644511149
transform 1 0 13708 0 -1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_179_149
timestamp 1644511149
transform 1 0 14812 0 -1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_179_161
timestamp 1644511149
transform 1 0 15916 0 -1 100096
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_179_167
timestamp 1644511149
transform 1 0 16468 0 -1 100096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_179_169
timestamp 1644511149
transform 1 0 16652 0 -1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_179_181
timestamp 1644511149
transform 1 0 17756 0 -1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_179_193
timestamp 1644511149
transform 1 0 18860 0 -1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_179_205
timestamp 1644511149
transform 1 0 19964 0 -1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_179_217
timestamp 1644511149
transform 1 0 21068 0 -1 100096
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_179_223
timestamp 1644511149
transform 1 0 21620 0 -1 100096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_179_225
timestamp 1644511149
transform 1 0 21804 0 -1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_179_237
timestamp 1644511149
transform 1 0 22908 0 -1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_179_249
timestamp 1644511149
transform 1 0 24012 0 -1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_179_261
timestamp 1644511149
transform 1 0 25116 0 -1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_179_273
timestamp 1644511149
transform 1 0 26220 0 -1 100096
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_179_279
timestamp 1644511149
transform 1 0 26772 0 -1 100096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_179_281
timestamp 1644511149
transform 1 0 26956 0 -1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_179_293
timestamp 1644511149
transform 1 0 28060 0 -1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_179_305
timestamp 1644511149
transform 1 0 29164 0 -1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_179_317
timestamp 1644511149
transform 1 0 30268 0 -1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_179_329
timestamp 1644511149
transform 1 0 31372 0 -1 100096
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_179_335
timestamp 1644511149
transform 1 0 31924 0 -1 100096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_179_337
timestamp 1644511149
transform 1 0 32108 0 -1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_179_349
timestamp 1644511149
transform 1 0 33212 0 -1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_179_361
timestamp 1644511149
transform 1 0 34316 0 -1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_179_373
timestamp 1644511149
transform 1 0 35420 0 -1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_179_385
timestamp 1644511149
transform 1 0 36524 0 -1 100096
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_179_391
timestamp 1644511149
transform 1 0 37076 0 -1 100096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_179_393
timestamp 1644511149
transform 1 0 37260 0 -1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_179_405
timestamp 1644511149
transform 1 0 38364 0 -1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_179_417
timestamp 1644511149
transform 1 0 39468 0 -1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_179_429
timestamp 1644511149
transform 1 0 40572 0 -1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_179_441
timestamp 1644511149
transform 1 0 41676 0 -1 100096
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_179_447
timestamp 1644511149
transform 1 0 42228 0 -1 100096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_179_449
timestamp 1644511149
transform 1 0 42412 0 -1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_179_461
timestamp 1644511149
transform 1 0 43516 0 -1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_179_473
timestamp 1644511149
transform 1 0 44620 0 -1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_179_485
timestamp 1644511149
transform 1 0 45724 0 -1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_179_497
timestamp 1644511149
transform 1 0 46828 0 -1 100096
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_179_503
timestamp 1644511149
transform 1 0 47380 0 -1 100096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_179_505
timestamp 1644511149
transform 1 0 47564 0 -1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_179_517
timestamp 1644511149
transform 1 0 48668 0 -1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_179_529
timestamp 1644511149
transform 1 0 49772 0 -1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_179_541
timestamp 1644511149
transform 1 0 50876 0 -1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_179_553
timestamp 1644511149
transform 1 0 51980 0 -1 100096
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_179_559
timestamp 1644511149
transform 1 0 52532 0 -1 100096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_179_561
timestamp 1644511149
transform 1 0 52716 0 -1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_179_573
timestamp 1644511149
transform 1 0 53820 0 -1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_179_585
timestamp 1644511149
transform 1 0 54924 0 -1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_179_597
timestamp 1644511149
transform 1 0 56028 0 -1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_179_609
timestamp 1644511149
transform 1 0 57132 0 -1 100096
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_179_615
timestamp 1644511149
transform 1 0 57684 0 -1 100096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_179_617
timestamp 1644511149
transform 1 0 57868 0 -1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_179_629
timestamp 1644511149
transform 1 0 58972 0 -1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_179_641
timestamp 1644511149
transform 1 0 60076 0 -1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_179_653
timestamp 1644511149
transform 1 0 61180 0 -1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_179_665
timestamp 1644511149
transform 1 0 62284 0 -1 100096
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_179_671
timestamp 1644511149
transform 1 0 62836 0 -1 100096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_179_673
timestamp 1644511149
transform 1 0 63020 0 -1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_179_685
timestamp 1644511149
transform 1 0 64124 0 -1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_179_697
timestamp 1644511149
transform 1 0 65228 0 -1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_179_709
timestamp 1644511149
transform 1 0 66332 0 -1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_179_721
timestamp 1644511149
transform 1 0 67436 0 -1 100096
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_179_727
timestamp 1644511149
transform 1 0 67988 0 -1 100096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_179_729
timestamp 1644511149
transform 1 0 68172 0 -1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_179_741
timestamp 1644511149
transform 1 0 69276 0 -1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_179_753
timestamp 1644511149
transform 1 0 70380 0 -1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_179_765
timestamp 1644511149
transform 1 0 71484 0 -1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_179_777
timestamp 1644511149
transform 1 0 72588 0 -1 100096
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_179_783
timestamp 1644511149
transform 1 0 73140 0 -1 100096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_179_785
timestamp 1644511149
transform 1 0 73324 0 -1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_179_797
timestamp 1644511149
transform 1 0 74428 0 -1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_179_809
timestamp 1644511149
transform 1 0 75532 0 -1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_179_821
timestamp 1644511149
transform 1 0 76636 0 -1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_179_833
timestamp 1644511149
transform 1 0 77740 0 -1 100096
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_179_839
timestamp 1644511149
transform 1 0 78292 0 -1 100096
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_179_841
timestamp 1644511149
transform 1 0 78476 0 -1 100096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_180_3
timestamp 1644511149
transform 1 0 1380 0 1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_180_15
timestamp 1644511149
transform 1 0 2484 0 1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_180_27
timestamp 1644511149
transform 1 0 3588 0 1 100096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_180_29
timestamp 1644511149
transform 1 0 3772 0 1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_180_41
timestamp 1644511149
transform 1 0 4876 0 1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_180_53
timestamp 1644511149
transform 1 0 5980 0 1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_180_65
timestamp 1644511149
transform 1 0 7084 0 1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_180_77
timestamp 1644511149
transform 1 0 8188 0 1 100096
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_180_83
timestamp 1644511149
transform 1 0 8740 0 1 100096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_180_85
timestamp 1644511149
transform 1 0 8924 0 1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_180_97
timestamp 1644511149
transform 1 0 10028 0 1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_180_109
timestamp 1644511149
transform 1 0 11132 0 1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_180_121
timestamp 1644511149
transform 1 0 12236 0 1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_180_133
timestamp 1644511149
transform 1 0 13340 0 1 100096
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_180_139
timestamp 1644511149
transform 1 0 13892 0 1 100096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_180_141
timestamp 1644511149
transform 1 0 14076 0 1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_180_153
timestamp 1644511149
transform 1 0 15180 0 1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_180_165
timestamp 1644511149
transform 1 0 16284 0 1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_180_177
timestamp 1644511149
transform 1 0 17388 0 1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_180_189
timestamp 1644511149
transform 1 0 18492 0 1 100096
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_180_195
timestamp 1644511149
transform 1 0 19044 0 1 100096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_180_197
timestamp 1644511149
transform 1 0 19228 0 1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_180_209
timestamp 1644511149
transform 1 0 20332 0 1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_180_221
timestamp 1644511149
transform 1 0 21436 0 1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_180_233
timestamp 1644511149
transform 1 0 22540 0 1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_180_245
timestamp 1644511149
transform 1 0 23644 0 1 100096
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_180_251
timestamp 1644511149
transform 1 0 24196 0 1 100096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_180_253
timestamp 1644511149
transform 1 0 24380 0 1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_180_265
timestamp 1644511149
transform 1 0 25484 0 1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_180_277
timestamp 1644511149
transform 1 0 26588 0 1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_180_289
timestamp 1644511149
transform 1 0 27692 0 1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_180_301
timestamp 1644511149
transform 1 0 28796 0 1 100096
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_180_307
timestamp 1644511149
transform 1 0 29348 0 1 100096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_180_309
timestamp 1644511149
transform 1 0 29532 0 1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_180_321
timestamp 1644511149
transform 1 0 30636 0 1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_180_333
timestamp 1644511149
transform 1 0 31740 0 1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_180_345
timestamp 1644511149
transform 1 0 32844 0 1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_180_357
timestamp 1644511149
transform 1 0 33948 0 1 100096
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_180_363
timestamp 1644511149
transform 1 0 34500 0 1 100096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_180_365
timestamp 1644511149
transform 1 0 34684 0 1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_180_377
timestamp 1644511149
transform 1 0 35788 0 1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_180_389
timestamp 1644511149
transform 1 0 36892 0 1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_180_401
timestamp 1644511149
transform 1 0 37996 0 1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_180_413
timestamp 1644511149
transform 1 0 39100 0 1 100096
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_180_419
timestamp 1644511149
transform 1 0 39652 0 1 100096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_180_421
timestamp 1644511149
transform 1 0 39836 0 1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_180_433
timestamp 1644511149
transform 1 0 40940 0 1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_180_445
timestamp 1644511149
transform 1 0 42044 0 1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_180_457
timestamp 1644511149
transform 1 0 43148 0 1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_180_469
timestamp 1644511149
transform 1 0 44252 0 1 100096
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_180_475
timestamp 1644511149
transform 1 0 44804 0 1 100096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_180_477
timestamp 1644511149
transform 1 0 44988 0 1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_180_489
timestamp 1644511149
transform 1 0 46092 0 1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_180_501
timestamp 1644511149
transform 1 0 47196 0 1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_180_513
timestamp 1644511149
transform 1 0 48300 0 1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_180_525
timestamp 1644511149
transform 1 0 49404 0 1 100096
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_180_531
timestamp 1644511149
transform 1 0 49956 0 1 100096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_180_533
timestamp 1644511149
transform 1 0 50140 0 1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_180_545
timestamp 1644511149
transform 1 0 51244 0 1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_180_557
timestamp 1644511149
transform 1 0 52348 0 1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_180_569
timestamp 1644511149
transform 1 0 53452 0 1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_180_581
timestamp 1644511149
transform 1 0 54556 0 1 100096
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_180_587
timestamp 1644511149
transform 1 0 55108 0 1 100096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_180_589
timestamp 1644511149
transform 1 0 55292 0 1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_180_601
timestamp 1644511149
transform 1 0 56396 0 1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_180_613
timestamp 1644511149
transform 1 0 57500 0 1 100096
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_180_621
timestamp 1644511149
transform 1 0 58236 0 1 100096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_180_627
timestamp 1644511149
transform 1 0 58788 0 1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_180_639
timestamp 1644511149
transform 1 0 59892 0 1 100096
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_180_643
timestamp 1644511149
transform 1 0 60260 0 1 100096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_180_645
timestamp 1644511149
transform 1 0 60444 0 1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_180_657
timestamp 1644511149
transform 1 0 61548 0 1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_180_669
timestamp 1644511149
transform 1 0 62652 0 1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_180_681
timestamp 1644511149
transform 1 0 63756 0 1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_180_693
timestamp 1644511149
transform 1 0 64860 0 1 100096
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_180_699
timestamp 1644511149
transform 1 0 65412 0 1 100096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_180_701
timestamp 1644511149
transform 1 0 65596 0 1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_180_713
timestamp 1644511149
transform 1 0 66700 0 1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_180_725
timestamp 1644511149
transform 1 0 67804 0 1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_180_737
timestamp 1644511149
transform 1 0 68908 0 1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_180_749
timestamp 1644511149
transform 1 0 70012 0 1 100096
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_180_755
timestamp 1644511149
transform 1 0 70564 0 1 100096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_180_757
timestamp 1644511149
transform 1 0 70748 0 1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_180_769
timestamp 1644511149
transform 1 0 71852 0 1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_180_781
timestamp 1644511149
transform 1 0 72956 0 1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_180_793
timestamp 1644511149
transform 1 0 74060 0 1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_180_805
timestamp 1644511149
transform 1 0 75164 0 1 100096
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_180_811
timestamp 1644511149
transform 1 0 75716 0 1 100096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_180_813
timestamp 1644511149
transform 1 0 75900 0 1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_180_825
timestamp 1644511149
transform 1 0 77004 0 1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_180_837
timestamp 1644511149
transform 1 0 78108 0 1 100096
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_180_841
timestamp 1644511149
transform 1 0 78476 0 1 100096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_181_3
timestamp 1644511149
transform 1 0 1380 0 -1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_181_15
timestamp 1644511149
transform 1 0 2484 0 -1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_181_27
timestamp 1644511149
transform 1 0 3588 0 -1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_181_39
timestamp 1644511149
transform 1 0 4692 0 -1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_181_51
timestamp 1644511149
transform 1 0 5796 0 -1 101184
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_181_55
timestamp 1644511149
transform 1 0 6164 0 -1 101184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_181_57
timestamp 1644511149
transform 1 0 6348 0 -1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_181_69
timestamp 1644511149
transform 1 0 7452 0 -1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_181_81
timestamp 1644511149
transform 1 0 8556 0 -1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_181_93
timestamp 1644511149
transform 1 0 9660 0 -1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_181_105
timestamp 1644511149
transform 1 0 10764 0 -1 101184
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_181_111
timestamp 1644511149
transform 1 0 11316 0 -1 101184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_181_113
timestamp 1644511149
transform 1 0 11500 0 -1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_181_125
timestamp 1644511149
transform 1 0 12604 0 -1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_181_137
timestamp 1644511149
transform 1 0 13708 0 -1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_181_149
timestamp 1644511149
transform 1 0 14812 0 -1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_181_161
timestamp 1644511149
transform 1 0 15916 0 -1 101184
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_181_167
timestamp 1644511149
transform 1 0 16468 0 -1 101184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_181_169
timestamp 1644511149
transform 1 0 16652 0 -1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_181_181
timestamp 1644511149
transform 1 0 17756 0 -1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_181_193
timestamp 1644511149
transform 1 0 18860 0 -1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_181_205
timestamp 1644511149
transform 1 0 19964 0 -1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_181_217
timestamp 1644511149
transform 1 0 21068 0 -1 101184
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_181_223
timestamp 1644511149
transform 1 0 21620 0 -1 101184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_181_225
timestamp 1644511149
transform 1 0 21804 0 -1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_181_237
timestamp 1644511149
transform 1 0 22908 0 -1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_181_249
timestamp 1644511149
transform 1 0 24012 0 -1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_181_261
timestamp 1644511149
transform 1 0 25116 0 -1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_181_273
timestamp 1644511149
transform 1 0 26220 0 -1 101184
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_181_279
timestamp 1644511149
transform 1 0 26772 0 -1 101184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_181_281
timestamp 1644511149
transform 1 0 26956 0 -1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_181_293
timestamp 1644511149
transform 1 0 28060 0 -1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_181_305
timestamp 1644511149
transform 1 0 29164 0 -1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_181_317
timestamp 1644511149
transform 1 0 30268 0 -1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_181_329
timestamp 1644511149
transform 1 0 31372 0 -1 101184
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_181_335
timestamp 1644511149
transform 1 0 31924 0 -1 101184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_181_337
timestamp 1644511149
transform 1 0 32108 0 -1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_181_349
timestamp 1644511149
transform 1 0 33212 0 -1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_181_361
timestamp 1644511149
transform 1 0 34316 0 -1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_181_373
timestamp 1644511149
transform 1 0 35420 0 -1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_181_385
timestamp 1644511149
transform 1 0 36524 0 -1 101184
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_181_391
timestamp 1644511149
transform 1 0 37076 0 -1 101184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_181_393
timestamp 1644511149
transform 1 0 37260 0 -1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_181_405
timestamp 1644511149
transform 1 0 38364 0 -1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_181_417
timestamp 1644511149
transform 1 0 39468 0 -1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_181_429
timestamp 1644511149
transform 1 0 40572 0 -1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_181_441
timestamp 1644511149
transform 1 0 41676 0 -1 101184
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_181_447
timestamp 1644511149
transform 1 0 42228 0 -1 101184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_181_449
timestamp 1644511149
transform 1 0 42412 0 -1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_181_461
timestamp 1644511149
transform 1 0 43516 0 -1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_181_473
timestamp 1644511149
transform 1 0 44620 0 -1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_181_485
timestamp 1644511149
transform 1 0 45724 0 -1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_181_497
timestamp 1644511149
transform 1 0 46828 0 -1 101184
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_181_503
timestamp 1644511149
transform 1 0 47380 0 -1 101184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_181_505
timestamp 1644511149
transform 1 0 47564 0 -1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_181_517
timestamp 1644511149
transform 1 0 48668 0 -1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_181_529
timestamp 1644511149
transform 1 0 49772 0 -1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_181_541
timestamp 1644511149
transform 1 0 50876 0 -1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_181_553
timestamp 1644511149
transform 1 0 51980 0 -1 101184
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_181_559
timestamp 1644511149
transform 1 0 52532 0 -1 101184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_181_561
timestamp 1644511149
transform 1 0 52716 0 -1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_181_573
timestamp 1644511149
transform 1 0 53820 0 -1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_181_585
timestamp 1644511149
transform 1 0 54924 0 -1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_181_597
timestamp 1644511149
transform 1 0 56028 0 -1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_181_609
timestamp 1644511149
transform 1 0 57132 0 -1 101184
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_181_615
timestamp 1644511149
transform 1 0 57684 0 -1 101184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_181_617
timestamp 1644511149
transform 1 0 57868 0 -1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_181_629
timestamp 1644511149
transform 1 0 58972 0 -1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_181_641
timestamp 1644511149
transform 1 0 60076 0 -1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_181_653
timestamp 1644511149
transform 1 0 61180 0 -1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_181_665
timestamp 1644511149
transform 1 0 62284 0 -1 101184
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_181_671
timestamp 1644511149
transform 1 0 62836 0 -1 101184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_181_673
timestamp 1644511149
transform 1 0 63020 0 -1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_181_685
timestamp 1644511149
transform 1 0 64124 0 -1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_181_697
timestamp 1644511149
transform 1 0 65228 0 -1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_181_709
timestamp 1644511149
transform 1 0 66332 0 -1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_181_721
timestamp 1644511149
transform 1 0 67436 0 -1 101184
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_181_727
timestamp 1644511149
transform 1 0 67988 0 -1 101184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_181_729
timestamp 1644511149
transform 1 0 68172 0 -1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_181_741
timestamp 1644511149
transform 1 0 69276 0 -1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_181_753
timestamp 1644511149
transform 1 0 70380 0 -1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_181_765
timestamp 1644511149
transform 1 0 71484 0 -1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_181_777
timestamp 1644511149
transform 1 0 72588 0 -1 101184
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_181_783
timestamp 1644511149
transform 1 0 73140 0 -1 101184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_181_785
timestamp 1644511149
transform 1 0 73324 0 -1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_181_797
timestamp 1644511149
transform 1 0 74428 0 -1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_181_809
timestamp 1644511149
transform 1 0 75532 0 -1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_181_821
timestamp 1644511149
transform 1 0 76636 0 -1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_181_833
timestamp 1644511149
transform 1 0 77740 0 -1 101184
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_181_839
timestamp 1644511149
transform 1 0 78292 0 -1 101184
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_181_841
timestamp 1644511149
transform 1 0 78476 0 -1 101184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_182_7
timestamp 1644511149
transform 1 0 1748 0 1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_182_19
timestamp 1644511149
transform 1 0 2852 0 1 101184
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_182_27
timestamp 1644511149
transform 1 0 3588 0 1 101184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_182_29
timestamp 1644511149
transform 1 0 3772 0 1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_182_41
timestamp 1644511149
transform 1 0 4876 0 1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_182_53
timestamp 1644511149
transform 1 0 5980 0 1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_182_65
timestamp 1644511149
transform 1 0 7084 0 1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_182_77
timestamp 1644511149
transform 1 0 8188 0 1 101184
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_182_83
timestamp 1644511149
transform 1 0 8740 0 1 101184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_182_85
timestamp 1644511149
transform 1 0 8924 0 1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_182_97
timestamp 1644511149
transform 1 0 10028 0 1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_182_109
timestamp 1644511149
transform 1 0 11132 0 1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_182_121
timestamp 1644511149
transform 1 0 12236 0 1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_182_133
timestamp 1644511149
transform 1 0 13340 0 1 101184
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_182_139
timestamp 1644511149
transform 1 0 13892 0 1 101184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_182_141
timestamp 1644511149
transform 1 0 14076 0 1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_182_153
timestamp 1644511149
transform 1 0 15180 0 1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_182_165
timestamp 1644511149
transform 1 0 16284 0 1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_182_177
timestamp 1644511149
transform 1 0 17388 0 1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_182_189
timestamp 1644511149
transform 1 0 18492 0 1 101184
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_182_195
timestamp 1644511149
transform 1 0 19044 0 1 101184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_182_197
timestamp 1644511149
transform 1 0 19228 0 1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_182_209
timestamp 1644511149
transform 1 0 20332 0 1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_182_221
timestamp 1644511149
transform 1 0 21436 0 1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_182_233
timestamp 1644511149
transform 1 0 22540 0 1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_182_245
timestamp 1644511149
transform 1 0 23644 0 1 101184
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_182_251
timestamp 1644511149
transform 1 0 24196 0 1 101184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_182_253
timestamp 1644511149
transform 1 0 24380 0 1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_182_265
timestamp 1644511149
transform 1 0 25484 0 1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_182_277
timestamp 1644511149
transform 1 0 26588 0 1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_182_289
timestamp 1644511149
transform 1 0 27692 0 1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_182_301
timestamp 1644511149
transform 1 0 28796 0 1 101184
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_182_307
timestamp 1644511149
transform 1 0 29348 0 1 101184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_182_309
timestamp 1644511149
transform 1 0 29532 0 1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_182_321
timestamp 1644511149
transform 1 0 30636 0 1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_182_333
timestamp 1644511149
transform 1 0 31740 0 1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_182_345
timestamp 1644511149
transform 1 0 32844 0 1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_182_357
timestamp 1644511149
transform 1 0 33948 0 1 101184
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_182_363
timestamp 1644511149
transform 1 0 34500 0 1 101184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_182_365
timestamp 1644511149
transform 1 0 34684 0 1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_182_377
timestamp 1644511149
transform 1 0 35788 0 1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_182_389
timestamp 1644511149
transform 1 0 36892 0 1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_182_401
timestamp 1644511149
transform 1 0 37996 0 1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_182_413
timestamp 1644511149
transform 1 0 39100 0 1 101184
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_182_419
timestamp 1644511149
transform 1 0 39652 0 1 101184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_182_421
timestamp 1644511149
transform 1 0 39836 0 1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_182_433
timestamp 1644511149
transform 1 0 40940 0 1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_182_445
timestamp 1644511149
transform 1 0 42044 0 1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_182_457
timestamp 1644511149
transform 1 0 43148 0 1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_182_469
timestamp 1644511149
transform 1 0 44252 0 1 101184
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_182_475
timestamp 1644511149
transform 1 0 44804 0 1 101184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_182_477
timestamp 1644511149
transform 1 0 44988 0 1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_182_489
timestamp 1644511149
transform 1 0 46092 0 1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_182_501
timestamp 1644511149
transform 1 0 47196 0 1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_182_513
timestamp 1644511149
transform 1 0 48300 0 1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_182_525
timestamp 1644511149
transform 1 0 49404 0 1 101184
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_182_531
timestamp 1644511149
transform 1 0 49956 0 1 101184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_182_533
timestamp 1644511149
transform 1 0 50140 0 1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_182_545
timestamp 1644511149
transform 1 0 51244 0 1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_182_557
timestamp 1644511149
transform 1 0 52348 0 1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_182_569
timestamp 1644511149
transform 1 0 53452 0 1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_182_581
timestamp 1644511149
transform 1 0 54556 0 1 101184
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_182_587
timestamp 1644511149
transform 1 0 55108 0 1 101184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_182_589
timestamp 1644511149
transform 1 0 55292 0 1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_182_601
timestamp 1644511149
transform 1 0 56396 0 1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_182_613
timestamp 1644511149
transform 1 0 57500 0 1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_182_625
timestamp 1644511149
transform 1 0 58604 0 1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_182_637
timestamp 1644511149
transform 1 0 59708 0 1 101184
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_182_643
timestamp 1644511149
transform 1 0 60260 0 1 101184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_182_645
timestamp 1644511149
transform 1 0 60444 0 1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_182_657
timestamp 1644511149
transform 1 0 61548 0 1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_182_669
timestamp 1644511149
transform 1 0 62652 0 1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_182_681
timestamp 1644511149
transform 1 0 63756 0 1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_182_693
timestamp 1644511149
transform 1 0 64860 0 1 101184
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_182_699
timestamp 1644511149
transform 1 0 65412 0 1 101184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_182_701
timestamp 1644511149
transform 1 0 65596 0 1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_182_713
timestamp 1644511149
transform 1 0 66700 0 1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_182_725
timestamp 1644511149
transform 1 0 67804 0 1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_182_737
timestamp 1644511149
transform 1 0 68908 0 1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_182_749
timestamp 1644511149
transform 1 0 70012 0 1 101184
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_182_755
timestamp 1644511149
transform 1 0 70564 0 1 101184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_182_757
timestamp 1644511149
transform 1 0 70748 0 1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_182_769
timestamp 1644511149
transform 1 0 71852 0 1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_182_781
timestamp 1644511149
transform 1 0 72956 0 1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_182_793
timestamp 1644511149
transform 1 0 74060 0 1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_182_805
timestamp 1644511149
transform 1 0 75164 0 1 101184
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_182_811
timestamp 1644511149
transform 1 0 75716 0 1 101184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_182_813
timestamp 1644511149
transform 1 0 75900 0 1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_182_825
timestamp 1644511149
transform 1 0 77004 0 1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_182_837
timestamp 1644511149
transform 1 0 78108 0 1 101184
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_182_841
timestamp 1644511149
transform 1 0 78476 0 1 101184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_183_3
timestamp 1644511149
transform 1 0 1380 0 -1 102272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_183_15
timestamp 1644511149
transform 1 0 2484 0 -1 102272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_183_27
timestamp 1644511149
transform 1 0 3588 0 -1 102272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_183_39
timestamp 1644511149
transform 1 0 4692 0 -1 102272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_183_51
timestamp 1644511149
transform 1 0 5796 0 -1 102272
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_183_55
timestamp 1644511149
transform 1 0 6164 0 -1 102272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_183_57
timestamp 1644511149
transform 1 0 6348 0 -1 102272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_183_69
timestamp 1644511149
transform 1 0 7452 0 -1 102272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_183_81
timestamp 1644511149
transform 1 0 8556 0 -1 102272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_183_93
timestamp 1644511149
transform 1 0 9660 0 -1 102272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_183_105
timestamp 1644511149
transform 1 0 10764 0 -1 102272
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_183_111
timestamp 1644511149
transform 1 0 11316 0 -1 102272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_183_113
timestamp 1644511149
transform 1 0 11500 0 -1 102272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_183_125
timestamp 1644511149
transform 1 0 12604 0 -1 102272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_183_137
timestamp 1644511149
transform 1 0 13708 0 -1 102272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_183_149
timestamp 1644511149
transform 1 0 14812 0 -1 102272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_183_161
timestamp 1644511149
transform 1 0 15916 0 -1 102272
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_183_167
timestamp 1644511149
transform 1 0 16468 0 -1 102272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_183_169
timestamp 1644511149
transform 1 0 16652 0 -1 102272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_183_181
timestamp 1644511149
transform 1 0 17756 0 -1 102272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_183_193
timestamp 1644511149
transform 1 0 18860 0 -1 102272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_183_205
timestamp 1644511149
transform 1 0 19964 0 -1 102272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_183_217
timestamp 1644511149
transform 1 0 21068 0 -1 102272
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_183_223
timestamp 1644511149
transform 1 0 21620 0 -1 102272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_183_225
timestamp 1644511149
transform 1 0 21804 0 -1 102272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_183_237
timestamp 1644511149
transform 1 0 22908 0 -1 102272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_183_249
timestamp 1644511149
transform 1 0 24012 0 -1 102272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_183_261
timestamp 1644511149
transform 1 0 25116 0 -1 102272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_183_273
timestamp 1644511149
transform 1 0 26220 0 -1 102272
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_183_279
timestamp 1644511149
transform 1 0 26772 0 -1 102272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_183_281
timestamp 1644511149
transform 1 0 26956 0 -1 102272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_183_293
timestamp 1644511149
transform 1 0 28060 0 -1 102272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_183_305
timestamp 1644511149
transform 1 0 29164 0 -1 102272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_183_317
timestamp 1644511149
transform 1 0 30268 0 -1 102272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_183_329
timestamp 1644511149
transform 1 0 31372 0 -1 102272
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_183_335
timestamp 1644511149
transform 1 0 31924 0 -1 102272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_183_337
timestamp 1644511149
transform 1 0 32108 0 -1 102272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_183_349
timestamp 1644511149
transform 1 0 33212 0 -1 102272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_183_361
timestamp 1644511149
transform 1 0 34316 0 -1 102272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_183_373
timestamp 1644511149
transform 1 0 35420 0 -1 102272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_183_385
timestamp 1644511149
transform 1 0 36524 0 -1 102272
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_183_391
timestamp 1644511149
transform 1 0 37076 0 -1 102272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_183_393
timestamp 1644511149
transform 1 0 37260 0 -1 102272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_183_405
timestamp 1644511149
transform 1 0 38364 0 -1 102272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_183_417
timestamp 1644511149
transform 1 0 39468 0 -1 102272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_183_429
timestamp 1644511149
transform 1 0 40572 0 -1 102272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_183_441
timestamp 1644511149
transform 1 0 41676 0 -1 102272
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_183_447
timestamp 1644511149
transform 1 0 42228 0 -1 102272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_183_449
timestamp 1644511149
transform 1 0 42412 0 -1 102272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_183_461
timestamp 1644511149
transform 1 0 43516 0 -1 102272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_183_473
timestamp 1644511149
transform 1 0 44620 0 -1 102272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_183_485
timestamp 1644511149
transform 1 0 45724 0 -1 102272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_183_497
timestamp 1644511149
transform 1 0 46828 0 -1 102272
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_183_503
timestamp 1644511149
transform 1 0 47380 0 -1 102272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_183_505
timestamp 1644511149
transform 1 0 47564 0 -1 102272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_183_517
timestamp 1644511149
transform 1 0 48668 0 -1 102272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_183_529
timestamp 1644511149
transform 1 0 49772 0 -1 102272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_183_541
timestamp 1644511149
transform 1 0 50876 0 -1 102272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_183_553
timestamp 1644511149
transform 1 0 51980 0 -1 102272
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_183_559
timestamp 1644511149
transform 1 0 52532 0 -1 102272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_183_561
timestamp 1644511149
transform 1 0 52716 0 -1 102272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_183_573
timestamp 1644511149
transform 1 0 53820 0 -1 102272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_183_585
timestamp 1644511149
transform 1 0 54924 0 -1 102272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_183_597
timestamp 1644511149
transform 1 0 56028 0 -1 102272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_183_609
timestamp 1644511149
transform 1 0 57132 0 -1 102272
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_183_615
timestamp 1644511149
transform 1 0 57684 0 -1 102272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_183_617
timestamp 1644511149
transform 1 0 57868 0 -1 102272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_183_629
timestamp 1644511149
transform 1 0 58972 0 -1 102272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_183_641
timestamp 1644511149
transform 1 0 60076 0 -1 102272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_183_653
timestamp 1644511149
transform 1 0 61180 0 -1 102272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_183_665
timestamp 1644511149
transform 1 0 62284 0 -1 102272
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_183_671
timestamp 1644511149
transform 1 0 62836 0 -1 102272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_183_673
timestamp 1644511149
transform 1 0 63020 0 -1 102272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_183_685
timestamp 1644511149
transform 1 0 64124 0 -1 102272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_183_697
timestamp 1644511149
transform 1 0 65228 0 -1 102272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_183_709
timestamp 1644511149
transform 1 0 66332 0 -1 102272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_183_721
timestamp 1644511149
transform 1 0 67436 0 -1 102272
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_183_727
timestamp 1644511149
transform 1 0 67988 0 -1 102272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_183_729
timestamp 1644511149
transform 1 0 68172 0 -1 102272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_183_741
timestamp 1644511149
transform 1 0 69276 0 -1 102272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_183_753
timestamp 1644511149
transform 1 0 70380 0 -1 102272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_183_765
timestamp 1644511149
transform 1 0 71484 0 -1 102272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_183_777
timestamp 1644511149
transform 1 0 72588 0 -1 102272
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_183_783
timestamp 1644511149
transform 1 0 73140 0 -1 102272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_183_785
timestamp 1644511149
transform 1 0 73324 0 -1 102272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_183_797
timestamp 1644511149
transform 1 0 74428 0 -1 102272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_183_809
timestamp 1644511149
transform 1 0 75532 0 -1 102272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_183_821
timestamp 1644511149
transform 1 0 76636 0 -1 102272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_183_833
timestamp 1644511149
transform 1 0 77740 0 -1 102272
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_183_839
timestamp 1644511149
transform 1 0 78292 0 -1 102272
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_183_841
timestamp 1644511149
transform 1 0 78476 0 -1 102272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_184_3
timestamp 1644511149
transform 1 0 1380 0 1 102272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_184_15
timestamp 1644511149
transform 1 0 2484 0 1 102272
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_184_27
timestamp 1644511149
transform 1 0 3588 0 1 102272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_184_29
timestamp 1644511149
transform 1 0 3772 0 1 102272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_184_41
timestamp 1644511149
transform 1 0 4876 0 1 102272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_184_53
timestamp 1644511149
transform 1 0 5980 0 1 102272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_184_65
timestamp 1644511149
transform 1 0 7084 0 1 102272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_184_77
timestamp 1644511149
transform 1 0 8188 0 1 102272
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_184_83
timestamp 1644511149
transform 1 0 8740 0 1 102272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_184_85
timestamp 1644511149
transform 1 0 8924 0 1 102272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_184_97
timestamp 1644511149
transform 1 0 10028 0 1 102272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_184_109
timestamp 1644511149
transform 1 0 11132 0 1 102272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_184_121
timestamp 1644511149
transform 1 0 12236 0 1 102272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_184_133
timestamp 1644511149
transform 1 0 13340 0 1 102272
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_184_139
timestamp 1644511149
transform 1 0 13892 0 1 102272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_184_141
timestamp 1644511149
transform 1 0 14076 0 1 102272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_184_153
timestamp 1644511149
transform 1 0 15180 0 1 102272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_184_165
timestamp 1644511149
transform 1 0 16284 0 1 102272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_184_177
timestamp 1644511149
transform 1 0 17388 0 1 102272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_184_189
timestamp 1644511149
transform 1 0 18492 0 1 102272
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_184_195
timestamp 1644511149
transform 1 0 19044 0 1 102272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_184_197
timestamp 1644511149
transform 1 0 19228 0 1 102272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_184_209
timestamp 1644511149
transform 1 0 20332 0 1 102272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_184_221
timestamp 1644511149
transform 1 0 21436 0 1 102272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_184_233
timestamp 1644511149
transform 1 0 22540 0 1 102272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_184_245
timestamp 1644511149
transform 1 0 23644 0 1 102272
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_184_251
timestamp 1644511149
transform 1 0 24196 0 1 102272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_184_253
timestamp 1644511149
transform 1 0 24380 0 1 102272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_184_265
timestamp 1644511149
transform 1 0 25484 0 1 102272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_184_277
timestamp 1644511149
transform 1 0 26588 0 1 102272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_184_289
timestamp 1644511149
transform 1 0 27692 0 1 102272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_184_301
timestamp 1644511149
transform 1 0 28796 0 1 102272
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_184_307
timestamp 1644511149
transform 1 0 29348 0 1 102272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_184_309
timestamp 1644511149
transform 1 0 29532 0 1 102272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_184_321
timestamp 1644511149
transform 1 0 30636 0 1 102272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_184_333
timestamp 1644511149
transform 1 0 31740 0 1 102272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_184_345
timestamp 1644511149
transform 1 0 32844 0 1 102272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_184_357
timestamp 1644511149
transform 1 0 33948 0 1 102272
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_184_363
timestamp 1644511149
transform 1 0 34500 0 1 102272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_184_365
timestamp 1644511149
transform 1 0 34684 0 1 102272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_184_377
timestamp 1644511149
transform 1 0 35788 0 1 102272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_184_389
timestamp 1644511149
transform 1 0 36892 0 1 102272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_184_401
timestamp 1644511149
transform 1 0 37996 0 1 102272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_184_413
timestamp 1644511149
transform 1 0 39100 0 1 102272
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_184_419
timestamp 1644511149
transform 1 0 39652 0 1 102272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_184_421
timestamp 1644511149
transform 1 0 39836 0 1 102272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_184_433
timestamp 1644511149
transform 1 0 40940 0 1 102272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_184_445
timestamp 1644511149
transform 1 0 42044 0 1 102272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_184_457
timestamp 1644511149
transform 1 0 43148 0 1 102272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_184_469
timestamp 1644511149
transform 1 0 44252 0 1 102272
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_184_475
timestamp 1644511149
transform 1 0 44804 0 1 102272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_184_477
timestamp 1644511149
transform 1 0 44988 0 1 102272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_184_489
timestamp 1644511149
transform 1 0 46092 0 1 102272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_184_501
timestamp 1644511149
transform 1 0 47196 0 1 102272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_184_513
timestamp 1644511149
transform 1 0 48300 0 1 102272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_184_525
timestamp 1644511149
transform 1 0 49404 0 1 102272
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_184_531
timestamp 1644511149
transform 1 0 49956 0 1 102272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_184_533
timestamp 1644511149
transform 1 0 50140 0 1 102272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_184_545
timestamp 1644511149
transform 1 0 51244 0 1 102272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_184_557
timestamp 1644511149
transform 1 0 52348 0 1 102272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_184_569
timestamp 1644511149
transform 1 0 53452 0 1 102272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_184_581
timestamp 1644511149
transform 1 0 54556 0 1 102272
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_184_587
timestamp 1644511149
transform 1 0 55108 0 1 102272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_184_589
timestamp 1644511149
transform 1 0 55292 0 1 102272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_184_601
timestamp 1644511149
transform 1 0 56396 0 1 102272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_184_613
timestamp 1644511149
transform 1 0 57500 0 1 102272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_184_625
timestamp 1644511149
transform 1 0 58604 0 1 102272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_184_637
timestamp 1644511149
transform 1 0 59708 0 1 102272
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_184_643
timestamp 1644511149
transform 1 0 60260 0 1 102272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_184_645
timestamp 1644511149
transform 1 0 60444 0 1 102272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_184_657
timestamp 1644511149
transform 1 0 61548 0 1 102272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_184_669
timestamp 1644511149
transform 1 0 62652 0 1 102272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_184_681
timestamp 1644511149
transform 1 0 63756 0 1 102272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_184_693
timestamp 1644511149
transform 1 0 64860 0 1 102272
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_184_699
timestamp 1644511149
transform 1 0 65412 0 1 102272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_184_701
timestamp 1644511149
transform 1 0 65596 0 1 102272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_184_713
timestamp 1644511149
transform 1 0 66700 0 1 102272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_184_725
timestamp 1644511149
transform 1 0 67804 0 1 102272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_184_737
timestamp 1644511149
transform 1 0 68908 0 1 102272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_184_749
timestamp 1644511149
transform 1 0 70012 0 1 102272
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_184_755
timestamp 1644511149
transform 1 0 70564 0 1 102272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_184_757
timestamp 1644511149
transform 1 0 70748 0 1 102272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_184_769
timestamp 1644511149
transform 1 0 71852 0 1 102272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_184_781
timestamp 1644511149
transform 1 0 72956 0 1 102272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_184_793
timestamp 1644511149
transform 1 0 74060 0 1 102272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_184_805
timestamp 1644511149
transform 1 0 75164 0 1 102272
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_184_811
timestamp 1644511149
transform 1 0 75716 0 1 102272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_184_813
timestamp 1644511149
transform 1 0 75900 0 1 102272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_184_825
timestamp 1644511149
transform 1 0 77004 0 1 102272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_184_837
timestamp 1644511149
transform 1 0 78108 0 1 102272
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_184_841
timestamp 1644511149
transform 1 0 78476 0 1 102272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_185_3
timestamp 1644511149
transform 1 0 1380 0 -1 103360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_185_15
timestamp 1644511149
transform 1 0 2484 0 -1 103360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_185_27
timestamp 1644511149
transform 1 0 3588 0 -1 103360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_185_39
timestamp 1644511149
transform 1 0 4692 0 -1 103360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_185_51
timestamp 1644511149
transform 1 0 5796 0 -1 103360
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_185_55
timestamp 1644511149
transform 1 0 6164 0 -1 103360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_185_57
timestamp 1644511149
transform 1 0 6348 0 -1 103360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_185_69
timestamp 1644511149
transform 1 0 7452 0 -1 103360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_185_81
timestamp 1644511149
transform 1 0 8556 0 -1 103360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_185_93
timestamp 1644511149
transform 1 0 9660 0 -1 103360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_185_105
timestamp 1644511149
transform 1 0 10764 0 -1 103360
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_185_111
timestamp 1644511149
transform 1 0 11316 0 -1 103360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_185_113
timestamp 1644511149
transform 1 0 11500 0 -1 103360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_185_125
timestamp 1644511149
transform 1 0 12604 0 -1 103360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_185_137
timestamp 1644511149
transform 1 0 13708 0 -1 103360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_185_149
timestamp 1644511149
transform 1 0 14812 0 -1 103360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_185_161
timestamp 1644511149
transform 1 0 15916 0 -1 103360
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_185_167
timestamp 1644511149
transform 1 0 16468 0 -1 103360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_185_169
timestamp 1644511149
transform 1 0 16652 0 -1 103360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_185_181
timestamp 1644511149
transform 1 0 17756 0 -1 103360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_185_193
timestamp 1644511149
transform 1 0 18860 0 -1 103360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_185_205
timestamp 1644511149
transform 1 0 19964 0 -1 103360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_185_217
timestamp 1644511149
transform 1 0 21068 0 -1 103360
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_185_223
timestamp 1644511149
transform 1 0 21620 0 -1 103360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_185_225
timestamp 1644511149
transform 1 0 21804 0 -1 103360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_185_237
timestamp 1644511149
transform 1 0 22908 0 -1 103360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_185_249
timestamp 1644511149
transform 1 0 24012 0 -1 103360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_185_261
timestamp 1644511149
transform 1 0 25116 0 -1 103360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_185_273
timestamp 1644511149
transform 1 0 26220 0 -1 103360
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_185_279
timestamp 1644511149
transform 1 0 26772 0 -1 103360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_185_281
timestamp 1644511149
transform 1 0 26956 0 -1 103360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_185_293
timestamp 1644511149
transform 1 0 28060 0 -1 103360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_185_305
timestamp 1644511149
transform 1 0 29164 0 -1 103360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_185_317
timestamp 1644511149
transform 1 0 30268 0 -1 103360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_185_329
timestamp 1644511149
transform 1 0 31372 0 -1 103360
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_185_335
timestamp 1644511149
transform 1 0 31924 0 -1 103360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_185_337
timestamp 1644511149
transform 1 0 32108 0 -1 103360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_185_349
timestamp 1644511149
transform 1 0 33212 0 -1 103360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_185_361
timestamp 1644511149
transform 1 0 34316 0 -1 103360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_185_373
timestamp 1644511149
transform 1 0 35420 0 -1 103360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_185_385
timestamp 1644511149
transform 1 0 36524 0 -1 103360
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_185_391
timestamp 1644511149
transform 1 0 37076 0 -1 103360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_185_393
timestamp 1644511149
transform 1 0 37260 0 -1 103360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_185_405
timestamp 1644511149
transform 1 0 38364 0 -1 103360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_185_417
timestamp 1644511149
transform 1 0 39468 0 -1 103360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_185_429
timestamp 1644511149
transform 1 0 40572 0 -1 103360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_185_441
timestamp 1644511149
transform 1 0 41676 0 -1 103360
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_185_447
timestamp 1644511149
transform 1 0 42228 0 -1 103360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_185_449
timestamp 1644511149
transform 1 0 42412 0 -1 103360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_185_461
timestamp 1644511149
transform 1 0 43516 0 -1 103360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_185_473
timestamp 1644511149
transform 1 0 44620 0 -1 103360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_185_485
timestamp 1644511149
transform 1 0 45724 0 -1 103360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_185_497
timestamp 1644511149
transform 1 0 46828 0 -1 103360
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_185_503
timestamp 1644511149
transform 1 0 47380 0 -1 103360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_185_505
timestamp 1644511149
transform 1 0 47564 0 -1 103360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_185_517
timestamp 1644511149
transform 1 0 48668 0 -1 103360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_185_529
timestamp 1644511149
transform 1 0 49772 0 -1 103360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_185_541
timestamp 1644511149
transform 1 0 50876 0 -1 103360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_185_553
timestamp 1644511149
transform 1 0 51980 0 -1 103360
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_185_559
timestamp 1644511149
transform 1 0 52532 0 -1 103360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_185_561
timestamp 1644511149
transform 1 0 52716 0 -1 103360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_185_573
timestamp 1644511149
transform 1 0 53820 0 -1 103360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_185_585
timestamp 1644511149
transform 1 0 54924 0 -1 103360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_185_597
timestamp 1644511149
transform 1 0 56028 0 -1 103360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_185_609
timestamp 1644511149
transform 1 0 57132 0 -1 103360
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_185_615
timestamp 1644511149
transform 1 0 57684 0 -1 103360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_185_617
timestamp 1644511149
transform 1 0 57868 0 -1 103360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_185_629
timestamp 1644511149
transform 1 0 58972 0 -1 103360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_185_641
timestamp 1644511149
transform 1 0 60076 0 -1 103360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_185_653
timestamp 1644511149
transform 1 0 61180 0 -1 103360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_185_665
timestamp 1644511149
transform 1 0 62284 0 -1 103360
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_185_671
timestamp 1644511149
transform 1 0 62836 0 -1 103360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_185_673
timestamp 1644511149
transform 1 0 63020 0 -1 103360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_185_685
timestamp 1644511149
transform 1 0 64124 0 -1 103360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_185_697
timestamp 1644511149
transform 1 0 65228 0 -1 103360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_185_709
timestamp 1644511149
transform 1 0 66332 0 -1 103360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_185_721
timestamp 1644511149
transform 1 0 67436 0 -1 103360
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_185_727
timestamp 1644511149
transform 1 0 67988 0 -1 103360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_185_729
timestamp 1644511149
transform 1 0 68172 0 -1 103360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_185_741
timestamp 1644511149
transform 1 0 69276 0 -1 103360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_185_753
timestamp 1644511149
transform 1 0 70380 0 -1 103360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_185_765
timestamp 1644511149
transform 1 0 71484 0 -1 103360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_185_777
timestamp 1644511149
transform 1 0 72588 0 -1 103360
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_185_783
timestamp 1644511149
transform 1 0 73140 0 -1 103360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_185_785
timestamp 1644511149
transform 1 0 73324 0 -1 103360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_185_797
timestamp 1644511149
transform 1 0 74428 0 -1 103360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_185_809
timestamp 1644511149
transform 1 0 75532 0 -1 103360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_185_821
timestamp 1644511149
transform 1 0 76636 0 -1 103360
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_185_827
timestamp 1644511149
transform 1 0 77188 0 -1 103360
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_185_830
timestamp 1644511149
transform 1 0 77464 0 -1 103360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_185_836
timestamp 1644511149
transform 1 0 78016 0 -1 103360
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_185_841
timestamp 1644511149
transform 1 0 78476 0 -1 103360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_186_3
timestamp 1644511149
transform 1 0 1380 0 1 103360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_186_15
timestamp 1644511149
transform 1 0 2484 0 1 103360
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_186_27
timestamp 1644511149
transform 1 0 3588 0 1 103360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_186_29
timestamp 1644511149
transform 1 0 3772 0 1 103360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_186_41
timestamp 1644511149
transform 1 0 4876 0 1 103360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_186_53
timestamp 1644511149
transform 1 0 5980 0 1 103360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_186_65
timestamp 1644511149
transform 1 0 7084 0 1 103360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_186_77
timestamp 1644511149
transform 1 0 8188 0 1 103360
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_186_83
timestamp 1644511149
transform 1 0 8740 0 1 103360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_186_85
timestamp 1644511149
transform 1 0 8924 0 1 103360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_186_97
timestamp 1644511149
transform 1 0 10028 0 1 103360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_186_109
timestamp 1644511149
transform 1 0 11132 0 1 103360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_186_121
timestamp 1644511149
transform 1 0 12236 0 1 103360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_186_133
timestamp 1644511149
transform 1 0 13340 0 1 103360
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_186_139
timestamp 1644511149
transform 1 0 13892 0 1 103360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_186_141
timestamp 1644511149
transform 1 0 14076 0 1 103360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_186_153
timestamp 1644511149
transform 1 0 15180 0 1 103360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_186_165
timestamp 1644511149
transform 1 0 16284 0 1 103360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_186_177
timestamp 1644511149
transform 1 0 17388 0 1 103360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_186_189
timestamp 1644511149
transform 1 0 18492 0 1 103360
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_186_195
timestamp 1644511149
transform 1 0 19044 0 1 103360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_186_197
timestamp 1644511149
transform 1 0 19228 0 1 103360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_186_209
timestamp 1644511149
transform 1 0 20332 0 1 103360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_186_221
timestamp 1644511149
transform 1 0 21436 0 1 103360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_186_233
timestamp 1644511149
transform 1 0 22540 0 1 103360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_186_245
timestamp 1644511149
transform 1 0 23644 0 1 103360
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_186_251
timestamp 1644511149
transform 1 0 24196 0 1 103360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_186_253
timestamp 1644511149
transform 1 0 24380 0 1 103360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_186_265
timestamp 1644511149
transform 1 0 25484 0 1 103360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_186_277
timestamp 1644511149
transform 1 0 26588 0 1 103360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_186_289
timestamp 1644511149
transform 1 0 27692 0 1 103360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_186_301
timestamp 1644511149
transform 1 0 28796 0 1 103360
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_186_307
timestamp 1644511149
transform 1 0 29348 0 1 103360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_186_309
timestamp 1644511149
transform 1 0 29532 0 1 103360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_186_321
timestamp 1644511149
transform 1 0 30636 0 1 103360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_186_333
timestamp 1644511149
transform 1 0 31740 0 1 103360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_186_345
timestamp 1644511149
transform 1 0 32844 0 1 103360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_186_357
timestamp 1644511149
transform 1 0 33948 0 1 103360
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_186_363
timestamp 1644511149
transform 1 0 34500 0 1 103360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_186_365
timestamp 1644511149
transform 1 0 34684 0 1 103360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_186_377
timestamp 1644511149
transform 1 0 35788 0 1 103360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_186_389
timestamp 1644511149
transform 1 0 36892 0 1 103360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_186_401
timestamp 1644511149
transform 1 0 37996 0 1 103360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_186_413
timestamp 1644511149
transform 1 0 39100 0 1 103360
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_186_419
timestamp 1644511149
transform 1 0 39652 0 1 103360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_186_421
timestamp 1644511149
transform 1 0 39836 0 1 103360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_186_433
timestamp 1644511149
transform 1 0 40940 0 1 103360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_186_445
timestamp 1644511149
transform 1 0 42044 0 1 103360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_186_457
timestamp 1644511149
transform 1 0 43148 0 1 103360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_186_469
timestamp 1644511149
transform 1 0 44252 0 1 103360
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_186_475
timestamp 1644511149
transform 1 0 44804 0 1 103360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_186_477
timestamp 1644511149
transform 1 0 44988 0 1 103360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_186_489
timestamp 1644511149
transform 1 0 46092 0 1 103360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_186_501
timestamp 1644511149
transform 1 0 47196 0 1 103360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_186_513
timestamp 1644511149
transform 1 0 48300 0 1 103360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_186_525
timestamp 1644511149
transform 1 0 49404 0 1 103360
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_186_531
timestamp 1644511149
transform 1 0 49956 0 1 103360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_186_533
timestamp 1644511149
transform 1 0 50140 0 1 103360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_186_545
timestamp 1644511149
transform 1 0 51244 0 1 103360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_186_557
timestamp 1644511149
transform 1 0 52348 0 1 103360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_186_569
timestamp 1644511149
transform 1 0 53452 0 1 103360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_186_581
timestamp 1644511149
transform 1 0 54556 0 1 103360
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_186_587
timestamp 1644511149
transform 1 0 55108 0 1 103360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_186_589
timestamp 1644511149
transform 1 0 55292 0 1 103360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_186_601
timestamp 1644511149
transform 1 0 56396 0 1 103360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_186_613
timestamp 1644511149
transform 1 0 57500 0 1 103360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_186_625
timestamp 1644511149
transform 1 0 58604 0 1 103360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_186_637
timestamp 1644511149
transform 1 0 59708 0 1 103360
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_186_643
timestamp 1644511149
transform 1 0 60260 0 1 103360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_186_645
timestamp 1644511149
transform 1 0 60444 0 1 103360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_186_657
timestamp 1644511149
transform 1 0 61548 0 1 103360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_186_669
timestamp 1644511149
transform 1 0 62652 0 1 103360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_186_681
timestamp 1644511149
transform 1 0 63756 0 1 103360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_186_693
timestamp 1644511149
transform 1 0 64860 0 1 103360
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_186_699
timestamp 1644511149
transform 1 0 65412 0 1 103360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_186_701
timestamp 1644511149
transform 1 0 65596 0 1 103360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_186_713
timestamp 1644511149
transform 1 0 66700 0 1 103360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_186_725
timestamp 1644511149
transform 1 0 67804 0 1 103360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_186_737
timestamp 1644511149
transform 1 0 68908 0 1 103360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_186_749
timestamp 1644511149
transform 1 0 70012 0 1 103360
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_186_755
timestamp 1644511149
transform 1 0 70564 0 1 103360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_186_757
timestamp 1644511149
transform 1 0 70748 0 1 103360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_186_769
timestamp 1644511149
transform 1 0 71852 0 1 103360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_186_781
timestamp 1644511149
transform 1 0 72956 0 1 103360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_186_793
timestamp 1644511149
transform 1 0 74060 0 1 103360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_186_805
timestamp 1644511149
transform 1 0 75164 0 1 103360
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_186_811
timestamp 1644511149
transform 1 0 75716 0 1 103360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_186_813
timestamp 1644511149
transform 1 0 75900 0 1 103360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_186_825
timestamp 1644511149
transform 1 0 77004 0 1 103360
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_186_833
timestamp 1644511149
transform 1 0 77740 0 1 103360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_186_837
timestamp 1644511149
transform 1 0 78108 0 1 103360
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_186_841
timestamp 1644511149
transform 1 0 78476 0 1 103360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_187_3
timestamp 1644511149
transform 1 0 1380 0 -1 104448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_187_15
timestamp 1644511149
transform 1 0 2484 0 -1 104448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_187_27
timestamp 1644511149
transform 1 0 3588 0 -1 104448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_187_39
timestamp 1644511149
transform 1 0 4692 0 -1 104448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_187_51
timestamp 1644511149
transform 1 0 5796 0 -1 104448
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_187_55
timestamp 1644511149
transform 1 0 6164 0 -1 104448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_187_57
timestamp 1644511149
transform 1 0 6348 0 -1 104448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_187_69
timestamp 1644511149
transform 1 0 7452 0 -1 104448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_187_81
timestamp 1644511149
transform 1 0 8556 0 -1 104448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_187_93
timestamp 1644511149
transform 1 0 9660 0 -1 104448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_187_105
timestamp 1644511149
transform 1 0 10764 0 -1 104448
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_187_111
timestamp 1644511149
transform 1 0 11316 0 -1 104448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_187_113
timestamp 1644511149
transform 1 0 11500 0 -1 104448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_187_125
timestamp 1644511149
transform 1 0 12604 0 -1 104448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_187_137
timestamp 1644511149
transform 1 0 13708 0 -1 104448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_187_149
timestamp 1644511149
transform 1 0 14812 0 -1 104448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_187_161
timestamp 1644511149
transform 1 0 15916 0 -1 104448
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_187_167
timestamp 1644511149
transform 1 0 16468 0 -1 104448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_187_169
timestamp 1644511149
transform 1 0 16652 0 -1 104448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_187_181
timestamp 1644511149
transform 1 0 17756 0 -1 104448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_187_193
timestamp 1644511149
transform 1 0 18860 0 -1 104448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_187_205
timestamp 1644511149
transform 1 0 19964 0 -1 104448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_187_217
timestamp 1644511149
transform 1 0 21068 0 -1 104448
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_187_223
timestamp 1644511149
transform 1 0 21620 0 -1 104448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_187_225
timestamp 1644511149
transform 1 0 21804 0 -1 104448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_187_237
timestamp 1644511149
transform 1 0 22908 0 -1 104448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_187_249
timestamp 1644511149
transform 1 0 24012 0 -1 104448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_187_261
timestamp 1644511149
transform 1 0 25116 0 -1 104448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_187_273
timestamp 1644511149
transform 1 0 26220 0 -1 104448
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_187_279
timestamp 1644511149
transform 1 0 26772 0 -1 104448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_187_281
timestamp 1644511149
transform 1 0 26956 0 -1 104448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_187_293
timestamp 1644511149
transform 1 0 28060 0 -1 104448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_187_305
timestamp 1644511149
transform 1 0 29164 0 -1 104448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_187_317
timestamp 1644511149
transform 1 0 30268 0 -1 104448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_187_329
timestamp 1644511149
transform 1 0 31372 0 -1 104448
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_187_335
timestamp 1644511149
transform 1 0 31924 0 -1 104448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_187_337
timestamp 1644511149
transform 1 0 32108 0 -1 104448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_187_349
timestamp 1644511149
transform 1 0 33212 0 -1 104448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_187_361
timestamp 1644511149
transform 1 0 34316 0 -1 104448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_187_373
timestamp 1644511149
transform 1 0 35420 0 -1 104448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_187_385
timestamp 1644511149
transform 1 0 36524 0 -1 104448
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_187_391
timestamp 1644511149
transform 1 0 37076 0 -1 104448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_187_393
timestamp 1644511149
transform 1 0 37260 0 -1 104448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_187_405
timestamp 1644511149
transform 1 0 38364 0 -1 104448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_187_417
timestamp 1644511149
transform 1 0 39468 0 -1 104448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_187_429
timestamp 1644511149
transform 1 0 40572 0 -1 104448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_187_441
timestamp 1644511149
transform 1 0 41676 0 -1 104448
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_187_447
timestamp 1644511149
transform 1 0 42228 0 -1 104448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_187_449
timestamp 1644511149
transform 1 0 42412 0 -1 104448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_187_461
timestamp 1644511149
transform 1 0 43516 0 -1 104448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_187_473
timestamp 1644511149
transform 1 0 44620 0 -1 104448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_187_485
timestamp 1644511149
transform 1 0 45724 0 -1 104448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_187_497
timestamp 1644511149
transform 1 0 46828 0 -1 104448
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_187_503
timestamp 1644511149
transform 1 0 47380 0 -1 104448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_187_505
timestamp 1644511149
transform 1 0 47564 0 -1 104448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_187_517
timestamp 1644511149
transform 1 0 48668 0 -1 104448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_187_529
timestamp 1644511149
transform 1 0 49772 0 -1 104448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_187_541
timestamp 1644511149
transform 1 0 50876 0 -1 104448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_187_553
timestamp 1644511149
transform 1 0 51980 0 -1 104448
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_187_559
timestamp 1644511149
transform 1 0 52532 0 -1 104448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_187_561
timestamp 1644511149
transform 1 0 52716 0 -1 104448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_187_573
timestamp 1644511149
transform 1 0 53820 0 -1 104448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_187_585
timestamp 1644511149
transform 1 0 54924 0 -1 104448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_187_597
timestamp 1644511149
transform 1 0 56028 0 -1 104448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_187_609
timestamp 1644511149
transform 1 0 57132 0 -1 104448
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_187_615
timestamp 1644511149
transform 1 0 57684 0 -1 104448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_187_617
timestamp 1644511149
transform 1 0 57868 0 -1 104448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_187_629
timestamp 1644511149
transform 1 0 58972 0 -1 104448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_187_641
timestamp 1644511149
transform 1 0 60076 0 -1 104448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_187_653
timestamp 1644511149
transform 1 0 61180 0 -1 104448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_187_665
timestamp 1644511149
transform 1 0 62284 0 -1 104448
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_187_671
timestamp 1644511149
transform 1 0 62836 0 -1 104448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_187_673
timestamp 1644511149
transform 1 0 63020 0 -1 104448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_187_685
timestamp 1644511149
transform 1 0 64124 0 -1 104448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_187_697
timestamp 1644511149
transform 1 0 65228 0 -1 104448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_187_709
timestamp 1644511149
transform 1 0 66332 0 -1 104448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_187_721
timestamp 1644511149
transform 1 0 67436 0 -1 104448
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_187_727
timestamp 1644511149
transform 1 0 67988 0 -1 104448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_187_729
timestamp 1644511149
transform 1 0 68172 0 -1 104448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_187_741
timestamp 1644511149
transform 1 0 69276 0 -1 104448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_187_753
timestamp 1644511149
transform 1 0 70380 0 -1 104448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_187_765
timestamp 1644511149
transform 1 0 71484 0 -1 104448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_187_777
timestamp 1644511149
transform 1 0 72588 0 -1 104448
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_187_783
timestamp 1644511149
transform 1 0 73140 0 -1 104448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_187_785
timestamp 1644511149
transform 1 0 73324 0 -1 104448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_187_797
timestamp 1644511149
transform 1 0 74428 0 -1 104448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_187_809
timestamp 1644511149
transform 1 0 75532 0 -1 104448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_187_821
timestamp 1644511149
transform 1 0 76636 0 -1 104448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_187_833
timestamp 1644511149
transform 1 0 77740 0 -1 104448
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_187_839
timestamp 1644511149
transform 1 0 78292 0 -1 104448
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_187_841
timestamp 1644511149
transform 1 0 78476 0 -1 104448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_188_3
timestamp 1644511149
transform 1 0 1380 0 1 104448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_188_15
timestamp 1644511149
transform 1 0 2484 0 1 104448
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_188_27
timestamp 1644511149
transform 1 0 3588 0 1 104448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_188_29
timestamp 1644511149
transform 1 0 3772 0 1 104448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_188_41
timestamp 1644511149
transform 1 0 4876 0 1 104448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_188_53
timestamp 1644511149
transform 1 0 5980 0 1 104448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_188_65
timestamp 1644511149
transform 1 0 7084 0 1 104448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_188_77
timestamp 1644511149
transform 1 0 8188 0 1 104448
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_188_83
timestamp 1644511149
transform 1 0 8740 0 1 104448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_188_85
timestamp 1644511149
transform 1 0 8924 0 1 104448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_188_97
timestamp 1644511149
transform 1 0 10028 0 1 104448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_188_109
timestamp 1644511149
transform 1 0 11132 0 1 104448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_188_121
timestamp 1644511149
transform 1 0 12236 0 1 104448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_188_133
timestamp 1644511149
transform 1 0 13340 0 1 104448
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_188_139
timestamp 1644511149
transform 1 0 13892 0 1 104448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_188_141
timestamp 1644511149
transform 1 0 14076 0 1 104448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_188_153
timestamp 1644511149
transform 1 0 15180 0 1 104448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_188_165
timestamp 1644511149
transform 1 0 16284 0 1 104448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_188_177
timestamp 1644511149
transform 1 0 17388 0 1 104448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_188_189
timestamp 1644511149
transform 1 0 18492 0 1 104448
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_188_195
timestamp 1644511149
transform 1 0 19044 0 1 104448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_188_197
timestamp 1644511149
transform 1 0 19228 0 1 104448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_188_209
timestamp 1644511149
transform 1 0 20332 0 1 104448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_188_221
timestamp 1644511149
transform 1 0 21436 0 1 104448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_188_233
timestamp 1644511149
transform 1 0 22540 0 1 104448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_188_245
timestamp 1644511149
transform 1 0 23644 0 1 104448
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_188_251
timestamp 1644511149
transform 1 0 24196 0 1 104448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_188_253
timestamp 1644511149
transform 1 0 24380 0 1 104448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_188_265
timestamp 1644511149
transform 1 0 25484 0 1 104448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_188_277
timestamp 1644511149
transform 1 0 26588 0 1 104448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_188_289
timestamp 1644511149
transform 1 0 27692 0 1 104448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_188_301
timestamp 1644511149
transform 1 0 28796 0 1 104448
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_188_307
timestamp 1644511149
transform 1 0 29348 0 1 104448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_188_309
timestamp 1644511149
transform 1 0 29532 0 1 104448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_188_321
timestamp 1644511149
transform 1 0 30636 0 1 104448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_188_333
timestamp 1644511149
transform 1 0 31740 0 1 104448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_188_345
timestamp 1644511149
transform 1 0 32844 0 1 104448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_188_357
timestamp 1644511149
transform 1 0 33948 0 1 104448
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_188_363
timestamp 1644511149
transform 1 0 34500 0 1 104448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_188_365
timestamp 1644511149
transform 1 0 34684 0 1 104448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_188_377
timestamp 1644511149
transform 1 0 35788 0 1 104448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_188_389
timestamp 1644511149
transform 1 0 36892 0 1 104448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_188_401
timestamp 1644511149
transform 1 0 37996 0 1 104448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_188_413
timestamp 1644511149
transform 1 0 39100 0 1 104448
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_188_419
timestamp 1644511149
transform 1 0 39652 0 1 104448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_188_421
timestamp 1644511149
transform 1 0 39836 0 1 104448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_188_433
timestamp 1644511149
transform 1 0 40940 0 1 104448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_188_445
timestamp 1644511149
transform 1 0 42044 0 1 104448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_188_457
timestamp 1644511149
transform 1 0 43148 0 1 104448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_188_469
timestamp 1644511149
transform 1 0 44252 0 1 104448
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_188_475
timestamp 1644511149
transform 1 0 44804 0 1 104448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_188_477
timestamp 1644511149
transform 1 0 44988 0 1 104448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_188_489
timestamp 1644511149
transform 1 0 46092 0 1 104448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_188_501
timestamp 1644511149
transform 1 0 47196 0 1 104448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_188_513
timestamp 1644511149
transform 1 0 48300 0 1 104448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_188_525
timestamp 1644511149
transform 1 0 49404 0 1 104448
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_188_531
timestamp 1644511149
transform 1 0 49956 0 1 104448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_188_533
timestamp 1644511149
transform 1 0 50140 0 1 104448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_188_545
timestamp 1644511149
transform 1 0 51244 0 1 104448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_188_557
timestamp 1644511149
transform 1 0 52348 0 1 104448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_188_569
timestamp 1644511149
transform 1 0 53452 0 1 104448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_188_581
timestamp 1644511149
transform 1 0 54556 0 1 104448
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_188_587
timestamp 1644511149
transform 1 0 55108 0 1 104448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_188_589
timestamp 1644511149
transform 1 0 55292 0 1 104448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_188_601
timestamp 1644511149
transform 1 0 56396 0 1 104448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_188_613
timestamp 1644511149
transform 1 0 57500 0 1 104448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_188_625
timestamp 1644511149
transform 1 0 58604 0 1 104448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_188_637
timestamp 1644511149
transform 1 0 59708 0 1 104448
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_188_643
timestamp 1644511149
transform 1 0 60260 0 1 104448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_188_645
timestamp 1644511149
transform 1 0 60444 0 1 104448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_188_657
timestamp 1644511149
transform 1 0 61548 0 1 104448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_188_669
timestamp 1644511149
transform 1 0 62652 0 1 104448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_188_681
timestamp 1644511149
transform 1 0 63756 0 1 104448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_188_693
timestamp 1644511149
transform 1 0 64860 0 1 104448
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_188_699
timestamp 1644511149
transform 1 0 65412 0 1 104448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_188_701
timestamp 1644511149
transform 1 0 65596 0 1 104448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_188_713
timestamp 1644511149
transform 1 0 66700 0 1 104448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_188_725
timestamp 1644511149
transform 1 0 67804 0 1 104448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_188_737
timestamp 1644511149
transform 1 0 68908 0 1 104448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_188_749
timestamp 1644511149
transform 1 0 70012 0 1 104448
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_188_755
timestamp 1644511149
transform 1 0 70564 0 1 104448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_188_757
timestamp 1644511149
transform 1 0 70748 0 1 104448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_188_769
timestamp 1644511149
transform 1 0 71852 0 1 104448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_188_781
timestamp 1644511149
transform 1 0 72956 0 1 104448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_188_793
timestamp 1644511149
transform 1 0 74060 0 1 104448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_188_805
timestamp 1644511149
transform 1 0 75164 0 1 104448
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_188_811
timestamp 1644511149
transform 1 0 75716 0 1 104448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_188_813
timestamp 1644511149
transform 1 0 75900 0 1 104448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_188_825
timestamp 1644511149
transform 1 0 77004 0 1 104448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_188_837
timestamp 1644511149
transform 1 0 78108 0 1 104448
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_188_841
timestamp 1644511149
transform 1 0 78476 0 1 104448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_189_3
timestamp 1644511149
transform 1 0 1380 0 -1 105536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_189_15
timestamp 1644511149
transform 1 0 2484 0 -1 105536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_189_27
timestamp 1644511149
transform 1 0 3588 0 -1 105536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_189_39
timestamp 1644511149
transform 1 0 4692 0 -1 105536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_189_51
timestamp 1644511149
transform 1 0 5796 0 -1 105536
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_189_55
timestamp 1644511149
transform 1 0 6164 0 -1 105536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_189_57
timestamp 1644511149
transform 1 0 6348 0 -1 105536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_189_69
timestamp 1644511149
transform 1 0 7452 0 -1 105536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_189_81
timestamp 1644511149
transform 1 0 8556 0 -1 105536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_189_93
timestamp 1644511149
transform 1 0 9660 0 -1 105536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_189_105
timestamp 1644511149
transform 1 0 10764 0 -1 105536
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_189_111
timestamp 1644511149
transform 1 0 11316 0 -1 105536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_189_113
timestamp 1644511149
transform 1 0 11500 0 -1 105536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_189_125
timestamp 1644511149
transform 1 0 12604 0 -1 105536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_189_137
timestamp 1644511149
transform 1 0 13708 0 -1 105536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_189_149
timestamp 1644511149
transform 1 0 14812 0 -1 105536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_189_161
timestamp 1644511149
transform 1 0 15916 0 -1 105536
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_189_167
timestamp 1644511149
transform 1 0 16468 0 -1 105536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_189_169
timestamp 1644511149
transform 1 0 16652 0 -1 105536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_189_181
timestamp 1644511149
transform 1 0 17756 0 -1 105536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_189_193
timestamp 1644511149
transform 1 0 18860 0 -1 105536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_189_205
timestamp 1644511149
transform 1 0 19964 0 -1 105536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_189_217
timestamp 1644511149
transform 1 0 21068 0 -1 105536
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_189_223
timestamp 1644511149
transform 1 0 21620 0 -1 105536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_189_225
timestamp 1644511149
transform 1 0 21804 0 -1 105536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_189_237
timestamp 1644511149
transform 1 0 22908 0 -1 105536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_189_249
timestamp 1644511149
transform 1 0 24012 0 -1 105536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_189_261
timestamp 1644511149
transform 1 0 25116 0 -1 105536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_189_273
timestamp 1644511149
transform 1 0 26220 0 -1 105536
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_189_279
timestamp 1644511149
transform 1 0 26772 0 -1 105536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_189_281
timestamp 1644511149
transform 1 0 26956 0 -1 105536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_189_293
timestamp 1644511149
transform 1 0 28060 0 -1 105536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_189_305
timestamp 1644511149
transform 1 0 29164 0 -1 105536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_189_317
timestamp 1644511149
transform 1 0 30268 0 -1 105536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_189_329
timestamp 1644511149
transform 1 0 31372 0 -1 105536
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_189_335
timestamp 1644511149
transform 1 0 31924 0 -1 105536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_189_337
timestamp 1644511149
transform 1 0 32108 0 -1 105536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_189_349
timestamp 1644511149
transform 1 0 33212 0 -1 105536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_189_361
timestamp 1644511149
transform 1 0 34316 0 -1 105536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_189_373
timestamp 1644511149
transform 1 0 35420 0 -1 105536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_189_385
timestamp 1644511149
transform 1 0 36524 0 -1 105536
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_189_391
timestamp 1644511149
transform 1 0 37076 0 -1 105536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_189_393
timestamp 1644511149
transform 1 0 37260 0 -1 105536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_189_405
timestamp 1644511149
transform 1 0 38364 0 -1 105536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_189_417
timestamp 1644511149
transform 1 0 39468 0 -1 105536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_189_429
timestamp 1644511149
transform 1 0 40572 0 -1 105536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_189_441
timestamp 1644511149
transform 1 0 41676 0 -1 105536
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_189_447
timestamp 1644511149
transform 1 0 42228 0 -1 105536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_189_449
timestamp 1644511149
transform 1 0 42412 0 -1 105536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_189_461
timestamp 1644511149
transform 1 0 43516 0 -1 105536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_189_473
timestamp 1644511149
transform 1 0 44620 0 -1 105536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_189_485
timestamp 1644511149
transform 1 0 45724 0 -1 105536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_189_497
timestamp 1644511149
transform 1 0 46828 0 -1 105536
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_189_503
timestamp 1644511149
transform 1 0 47380 0 -1 105536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_189_505
timestamp 1644511149
transform 1 0 47564 0 -1 105536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_189_517
timestamp 1644511149
transform 1 0 48668 0 -1 105536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_189_529
timestamp 1644511149
transform 1 0 49772 0 -1 105536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_189_541
timestamp 1644511149
transform 1 0 50876 0 -1 105536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_189_553
timestamp 1644511149
transform 1 0 51980 0 -1 105536
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_189_559
timestamp 1644511149
transform 1 0 52532 0 -1 105536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_189_561
timestamp 1644511149
transform 1 0 52716 0 -1 105536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_189_573
timestamp 1644511149
transform 1 0 53820 0 -1 105536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_189_585
timestamp 1644511149
transform 1 0 54924 0 -1 105536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_189_597
timestamp 1644511149
transform 1 0 56028 0 -1 105536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_189_609
timestamp 1644511149
transform 1 0 57132 0 -1 105536
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_189_615
timestamp 1644511149
transform 1 0 57684 0 -1 105536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_189_617
timestamp 1644511149
transform 1 0 57868 0 -1 105536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_189_629
timestamp 1644511149
transform 1 0 58972 0 -1 105536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_189_641
timestamp 1644511149
transform 1 0 60076 0 -1 105536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_189_653
timestamp 1644511149
transform 1 0 61180 0 -1 105536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_189_665
timestamp 1644511149
transform 1 0 62284 0 -1 105536
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_189_671
timestamp 1644511149
transform 1 0 62836 0 -1 105536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_189_673
timestamp 1644511149
transform 1 0 63020 0 -1 105536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_189_685
timestamp 1644511149
transform 1 0 64124 0 -1 105536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_189_697
timestamp 1644511149
transform 1 0 65228 0 -1 105536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_189_709
timestamp 1644511149
transform 1 0 66332 0 -1 105536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_189_721
timestamp 1644511149
transform 1 0 67436 0 -1 105536
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_189_727
timestamp 1644511149
transform 1 0 67988 0 -1 105536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_189_729
timestamp 1644511149
transform 1 0 68172 0 -1 105536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_189_741
timestamp 1644511149
transform 1 0 69276 0 -1 105536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_189_753
timestamp 1644511149
transform 1 0 70380 0 -1 105536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_189_765
timestamp 1644511149
transform 1 0 71484 0 -1 105536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_189_777
timestamp 1644511149
transform 1 0 72588 0 -1 105536
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_189_783
timestamp 1644511149
transform 1 0 73140 0 -1 105536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_189_785
timestamp 1644511149
transform 1 0 73324 0 -1 105536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_189_797
timestamp 1644511149
transform 1 0 74428 0 -1 105536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_189_809
timestamp 1644511149
transform 1 0 75532 0 -1 105536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_189_821
timestamp 1644511149
transform 1 0 76636 0 -1 105536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_189_833
timestamp 1644511149
transform 1 0 77740 0 -1 105536
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_189_839
timestamp 1644511149
transform 1 0 78292 0 -1 105536
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_189_841
timestamp 1644511149
transform 1 0 78476 0 -1 105536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_190_9
timestamp 1644511149
transform 1 0 1932 0 1 105536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_190_21
timestamp 1644511149
transform 1 0 3036 0 1 105536
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_190_27
timestamp 1644511149
transform 1 0 3588 0 1 105536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_190_29
timestamp 1644511149
transform 1 0 3772 0 1 105536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_190_41
timestamp 1644511149
transform 1 0 4876 0 1 105536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_190_53
timestamp 1644511149
transform 1 0 5980 0 1 105536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_190_65
timestamp 1644511149
transform 1 0 7084 0 1 105536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_190_77
timestamp 1644511149
transform 1 0 8188 0 1 105536
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_190_83
timestamp 1644511149
transform 1 0 8740 0 1 105536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_190_85
timestamp 1644511149
transform 1 0 8924 0 1 105536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_190_97
timestamp 1644511149
transform 1 0 10028 0 1 105536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_190_109
timestamp 1644511149
transform 1 0 11132 0 1 105536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_190_121
timestamp 1644511149
transform 1 0 12236 0 1 105536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_190_133
timestamp 1644511149
transform 1 0 13340 0 1 105536
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_190_139
timestamp 1644511149
transform 1 0 13892 0 1 105536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_190_141
timestamp 1644511149
transform 1 0 14076 0 1 105536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_190_153
timestamp 1644511149
transform 1 0 15180 0 1 105536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_190_165
timestamp 1644511149
transform 1 0 16284 0 1 105536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_190_177
timestamp 1644511149
transform 1 0 17388 0 1 105536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_190_189
timestamp 1644511149
transform 1 0 18492 0 1 105536
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_190_195
timestamp 1644511149
transform 1 0 19044 0 1 105536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_190_197
timestamp 1644511149
transform 1 0 19228 0 1 105536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_190_209
timestamp 1644511149
transform 1 0 20332 0 1 105536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_190_221
timestamp 1644511149
transform 1 0 21436 0 1 105536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_190_233
timestamp 1644511149
transform 1 0 22540 0 1 105536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_190_245
timestamp 1644511149
transform 1 0 23644 0 1 105536
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_190_251
timestamp 1644511149
transform 1 0 24196 0 1 105536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_190_253
timestamp 1644511149
transform 1 0 24380 0 1 105536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_190_265
timestamp 1644511149
transform 1 0 25484 0 1 105536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_190_277
timestamp 1644511149
transform 1 0 26588 0 1 105536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_190_289
timestamp 1644511149
transform 1 0 27692 0 1 105536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_190_301
timestamp 1644511149
transform 1 0 28796 0 1 105536
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_190_307
timestamp 1644511149
transform 1 0 29348 0 1 105536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_190_309
timestamp 1644511149
transform 1 0 29532 0 1 105536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_190_321
timestamp 1644511149
transform 1 0 30636 0 1 105536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_190_333
timestamp 1644511149
transform 1 0 31740 0 1 105536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_190_345
timestamp 1644511149
transform 1 0 32844 0 1 105536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_190_357
timestamp 1644511149
transform 1 0 33948 0 1 105536
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_190_363
timestamp 1644511149
transform 1 0 34500 0 1 105536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_190_365
timestamp 1644511149
transform 1 0 34684 0 1 105536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_190_377
timestamp 1644511149
transform 1 0 35788 0 1 105536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_190_389
timestamp 1644511149
transform 1 0 36892 0 1 105536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_190_401
timestamp 1644511149
transform 1 0 37996 0 1 105536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_190_413
timestamp 1644511149
transform 1 0 39100 0 1 105536
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_190_419
timestamp 1644511149
transform 1 0 39652 0 1 105536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_190_421
timestamp 1644511149
transform 1 0 39836 0 1 105536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_190_433
timestamp 1644511149
transform 1 0 40940 0 1 105536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_190_445
timestamp 1644511149
transform 1 0 42044 0 1 105536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_190_457
timestamp 1644511149
transform 1 0 43148 0 1 105536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_190_469
timestamp 1644511149
transform 1 0 44252 0 1 105536
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_190_475
timestamp 1644511149
transform 1 0 44804 0 1 105536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_190_477
timestamp 1644511149
transform 1 0 44988 0 1 105536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_190_489
timestamp 1644511149
transform 1 0 46092 0 1 105536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_190_501
timestamp 1644511149
transform 1 0 47196 0 1 105536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_190_513
timestamp 1644511149
transform 1 0 48300 0 1 105536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_190_525
timestamp 1644511149
transform 1 0 49404 0 1 105536
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_190_531
timestamp 1644511149
transform 1 0 49956 0 1 105536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_190_533
timestamp 1644511149
transform 1 0 50140 0 1 105536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_190_545
timestamp 1644511149
transform 1 0 51244 0 1 105536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_190_557
timestamp 1644511149
transform 1 0 52348 0 1 105536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_190_569
timestamp 1644511149
transform 1 0 53452 0 1 105536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_190_581
timestamp 1644511149
transform 1 0 54556 0 1 105536
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_190_587
timestamp 1644511149
transform 1 0 55108 0 1 105536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_190_589
timestamp 1644511149
transform 1 0 55292 0 1 105536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_190_601
timestamp 1644511149
transform 1 0 56396 0 1 105536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_190_613
timestamp 1644511149
transform 1 0 57500 0 1 105536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_190_625
timestamp 1644511149
transform 1 0 58604 0 1 105536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_190_637
timestamp 1644511149
transform 1 0 59708 0 1 105536
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_190_643
timestamp 1644511149
transform 1 0 60260 0 1 105536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_190_645
timestamp 1644511149
transform 1 0 60444 0 1 105536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_190_657
timestamp 1644511149
transform 1 0 61548 0 1 105536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_190_669
timestamp 1644511149
transform 1 0 62652 0 1 105536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_190_681
timestamp 1644511149
transform 1 0 63756 0 1 105536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_190_693
timestamp 1644511149
transform 1 0 64860 0 1 105536
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_190_699
timestamp 1644511149
transform 1 0 65412 0 1 105536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_190_701
timestamp 1644511149
transform 1 0 65596 0 1 105536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_190_713
timestamp 1644511149
transform 1 0 66700 0 1 105536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_190_725
timestamp 1644511149
transform 1 0 67804 0 1 105536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_190_737
timestamp 1644511149
transform 1 0 68908 0 1 105536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_190_749
timestamp 1644511149
transform 1 0 70012 0 1 105536
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_190_755
timestamp 1644511149
transform 1 0 70564 0 1 105536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_190_757
timestamp 1644511149
transform 1 0 70748 0 1 105536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_190_769
timestamp 1644511149
transform 1 0 71852 0 1 105536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_190_781
timestamp 1644511149
transform 1 0 72956 0 1 105536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_190_793
timestamp 1644511149
transform 1 0 74060 0 1 105536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_190_805
timestamp 1644511149
transform 1 0 75164 0 1 105536
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_190_811
timestamp 1644511149
transform 1 0 75716 0 1 105536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_190_813
timestamp 1644511149
transform 1 0 75900 0 1 105536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_190_825
timestamp 1644511149
transform 1 0 77004 0 1 105536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_190_837
timestamp 1644511149
transform 1 0 78108 0 1 105536
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_190_841
timestamp 1644511149
transform 1 0 78476 0 1 105536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_191_3
timestamp 1644511149
transform 1 0 1380 0 -1 106624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_191_15
timestamp 1644511149
transform 1 0 2484 0 -1 106624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_191_27
timestamp 1644511149
transform 1 0 3588 0 -1 106624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_191_39
timestamp 1644511149
transform 1 0 4692 0 -1 106624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_191_51
timestamp 1644511149
transform 1 0 5796 0 -1 106624
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_191_55
timestamp 1644511149
transform 1 0 6164 0 -1 106624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_191_57
timestamp 1644511149
transform 1 0 6348 0 -1 106624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_191_69
timestamp 1644511149
transform 1 0 7452 0 -1 106624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_191_81
timestamp 1644511149
transform 1 0 8556 0 -1 106624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_191_93
timestamp 1644511149
transform 1 0 9660 0 -1 106624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_191_105
timestamp 1644511149
transform 1 0 10764 0 -1 106624
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_191_111
timestamp 1644511149
transform 1 0 11316 0 -1 106624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_191_113
timestamp 1644511149
transform 1 0 11500 0 -1 106624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_191_125
timestamp 1644511149
transform 1 0 12604 0 -1 106624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_191_137
timestamp 1644511149
transform 1 0 13708 0 -1 106624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_191_149
timestamp 1644511149
transform 1 0 14812 0 -1 106624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_191_161
timestamp 1644511149
transform 1 0 15916 0 -1 106624
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_191_167
timestamp 1644511149
transform 1 0 16468 0 -1 106624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_191_169
timestamp 1644511149
transform 1 0 16652 0 -1 106624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_191_181
timestamp 1644511149
transform 1 0 17756 0 -1 106624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_191_193
timestamp 1644511149
transform 1 0 18860 0 -1 106624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_191_205
timestamp 1644511149
transform 1 0 19964 0 -1 106624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_191_217
timestamp 1644511149
transform 1 0 21068 0 -1 106624
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_191_223
timestamp 1644511149
transform 1 0 21620 0 -1 106624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_191_225
timestamp 1644511149
transform 1 0 21804 0 -1 106624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_191_237
timestamp 1644511149
transform 1 0 22908 0 -1 106624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_191_249
timestamp 1644511149
transform 1 0 24012 0 -1 106624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_191_261
timestamp 1644511149
transform 1 0 25116 0 -1 106624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_191_273
timestamp 1644511149
transform 1 0 26220 0 -1 106624
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_191_279
timestamp 1644511149
transform 1 0 26772 0 -1 106624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_191_281
timestamp 1644511149
transform 1 0 26956 0 -1 106624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_191_293
timestamp 1644511149
transform 1 0 28060 0 -1 106624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_191_305
timestamp 1644511149
transform 1 0 29164 0 -1 106624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_191_317
timestamp 1644511149
transform 1 0 30268 0 -1 106624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_191_329
timestamp 1644511149
transform 1 0 31372 0 -1 106624
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_191_335
timestamp 1644511149
transform 1 0 31924 0 -1 106624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_191_337
timestamp 1644511149
transform 1 0 32108 0 -1 106624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_191_349
timestamp 1644511149
transform 1 0 33212 0 -1 106624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_191_361
timestamp 1644511149
transform 1 0 34316 0 -1 106624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_191_373
timestamp 1644511149
transform 1 0 35420 0 -1 106624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_191_385
timestamp 1644511149
transform 1 0 36524 0 -1 106624
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_191_391
timestamp 1644511149
transform 1 0 37076 0 -1 106624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_191_393
timestamp 1644511149
transform 1 0 37260 0 -1 106624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_191_405
timestamp 1644511149
transform 1 0 38364 0 -1 106624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_191_417
timestamp 1644511149
transform 1 0 39468 0 -1 106624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_191_429
timestamp 1644511149
transform 1 0 40572 0 -1 106624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_191_441
timestamp 1644511149
transform 1 0 41676 0 -1 106624
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_191_447
timestamp 1644511149
transform 1 0 42228 0 -1 106624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_191_449
timestamp 1644511149
transform 1 0 42412 0 -1 106624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_191_461
timestamp 1644511149
transform 1 0 43516 0 -1 106624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_191_473
timestamp 1644511149
transform 1 0 44620 0 -1 106624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_191_485
timestamp 1644511149
transform 1 0 45724 0 -1 106624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_191_497
timestamp 1644511149
transform 1 0 46828 0 -1 106624
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_191_503
timestamp 1644511149
transform 1 0 47380 0 -1 106624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_191_505
timestamp 1644511149
transform 1 0 47564 0 -1 106624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_191_517
timestamp 1644511149
transform 1 0 48668 0 -1 106624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_191_529
timestamp 1644511149
transform 1 0 49772 0 -1 106624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_191_541
timestamp 1644511149
transform 1 0 50876 0 -1 106624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_191_553
timestamp 1644511149
transform 1 0 51980 0 -1 106624
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_191_559
timestamp 1644511149
transform 1 0 52532 0 -1 106624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_191_561
timestamp 1644511149
transform 1 0 52716 0 -1 106624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_191_573
timestamp 1644511149
transform 1 0 53820 0 -1 106624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_191_585
timestamp 1644511149
transform 1 0 54924 0 -1 106624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_191_597
timestamp 1644511149
transform 1 0 56028 0 -1 106624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_191_609
timestamp 1644511149
transform 1 0 57132 0 -1 106624
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_191_615
timestamp 1644511149
transform 1 0 57684 0 -1 106624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_191_617
timestamp 1644511149
transform 1 0 57868 0 -1 106624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_191_629
timestamp 1644511149
transform 1 0 58972 0 -1 106624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_191_641
timestamp 1644511149
transform 1 0 60076 0 -1 106624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_191_653
timestamp 1644511149
transform 1 0 61180 0 -1 106624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_191_665
timestamp 1644511149
transform 1 0 62284 0 -1 106624
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_191_671
timestamp 1644511149
transform 1 0 62836 0 -1 106624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_191_673
timestamp 1644511149
transform 1 0 63020 0 -1 106624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_191_685
timestamp 1644511149
transform 1 0 64124 0 -1 106624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_191_697
timestamp 1644511149
transform 1 0 65228 0 -1 106624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_191_709
timestamp 1644511149
transform 1 0 66332 0 -1 106624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_191_721
timestamp 1644511149
transform 1 0 67436 0 -1 106624
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_191_727
timestamp 1644511149
transform 1 0 67988 0 -1 106624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_191_729
timestamp 1644511149
transform 1 0 68172 0 -1 106624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_191_741
timestamp 1644511149
transform 1 0 69276 0 -1 106624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_191_753
timestamp 1644511149
transform 1 0 70380 0 -1 106624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_191_765
timestamp 1644511149
transform 1 0 71484 0 -1 106624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_191_777
timestamp 1644511149
transform 1 0 72588 0 -1 106624
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_191_783
timestamp 1644511149
transform 1 0 73140 0 -1 106624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_191_785
timestamp 1644511149
transform 1 0 73324 0 -1 106624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_191_797
timestamp 1644511149
transform 1 0 74428 0 -1 106624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_191_809
timestamp 1644511149
transform 1 0 75532 0 -1 106624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_191_821
timestamp 1644511149
transform 1 0 76636 0 -1 106624
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_191_829
timestamp 1644511149
transform 1 0 77372 0 -1 106624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_191_836
timestamp 1644511149
transform 1 0 78016 0 -1 106624
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_191_841
timestamp 1644511149
transform 1 0 78476 0 -1 106624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_192_3
timestamp 1644511149
transform 1 0 1380 0 1 106624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_192_15
timestamp 1644511149
transform 1 0 2484 0 1 106624
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_192_27
timestamp 1644511149
transform 1 0 3588 0 1 106624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_192_29
timestamp 1644511149
transform 1 0 3772 0 1 106624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_192_41
timestamp 1644511149
transform 1 0 4876 0 1 106624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_192_53
timestamp 1644511149
transform 1 0 5980 0 1 106624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_192_65
timestamp 1644511149
transform 1 0 7084 0 1 106624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_192_77
timestamp 1644511149
transform 1 0 8188 0 1 106624
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_192_83
timestamp 1644511149
transform 1 0 8740 0 1 106624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_192_85
timestamp 1644511149
transform 1 0 8924 0 1 106624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_192_97
timestamp 1644511149
transform 1 0 10028 0 1 106624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_192_109
timestamp 1644511149
transform 1 0 11132 0 1 106624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_192_121
timestamp 1644511149
transform 1 0 12236 0 1 106624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_192_133
timestamp 1644511149
transform 1 0 13340 0 1 106624
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_192_139
timestamp 1644511149
transform 1 0 13892 0 1 106624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_192_141
timestamp 1644511149
transform 1 0 14076 0 1 106624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_192_153
timestamp 1644511149
transform 1 0 15180 0 1 106624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_192_165
timestamp 1644511149
transform 1 0 16284 0 1 106624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_192_177
timestamp 1644511149
transform 1 0 17388 0 1 106624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_192_189
timestamp 1644511149
transform 1 0 18492 0 1 106624
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_192_195
timestamp 1644511149
transform 1 0 19044 0 1 106624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_192_197
timestamp 1644511149
transform 1 0 19228 0 1 106624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_192_209
timestamp 1644511149
transform 1 0 20332 0 1 106624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_192_221
timestamp 1644511149
transform 1 0 21436 0 1 106624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_192_233
timestamp 1644511149
transform 1 0 22540 0 1 106624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_192_245
timestamp 1644511149
transform 1 0 23644 0 1 106624
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_192_251
timestamp 1644511149
transform 1 0 24196 0 1 106624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_192_253
timestamp 1644511149
transform 1 0 24380 0 1 106624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_192_265
timestamp 1644511149
transform 1 0 25484 0 1 106624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_192_277
timestamp 1644511149
transform 1 0 26588 0 1 106624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_192_289
timestamp 1644511149
transform 1 0 27692 0 1 106624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_192_301
timestamp 1644511149
transform 1 0 28796 0 1 106624
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_192_307
timestamp 1644511149
transform 1 0 29348 0 1 106624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_192_309
timestamp 1644511149
transform 1 0 29532 0 1 106624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_192_321
timestamp 1644511149
transform 1 0 30636 0 1 106624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_192_333
timestamp 1644511149
transform 1 0 31740 0 1 106624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_192_345
timestamp 1644511149
transform 1 0 32844 0 1 106624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_192_357
timestamp 1644511149
transform 1 0 33948 0 1 106624
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_192_363
timestamp 1644511149
transform 1 0 34500 0 1 106624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_192_365
timestamp 1644511149
transform 1 0 34684 0 1 106624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_192_377
timestamp 1644511149
transform 1 0 35788 0 1 106624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_192_389
timestamp 1644511149
transform 1 0 36892 0 1 106624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_192_401
timestamp 1644511149
transform 1 0 37996 0 1 106624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_192_413
timestamp 1644511149
transform 1 0 39100 0 1 106624
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_192_419
timestamp 1644511149
transform 1 0 39652 0 1 106624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_192_421
timestamp 1644511149
transform 1 0 39836 0 1 106624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_192_433
timestamp 1644511149
transform 1 0 40940 0 1 106624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_192_445
timestamp 1644511149
transform 1 0 42044 0 1 106624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_192_457
timestamp 1644511149
transform 1 0 43148 0 1 106624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_192_469
timestamp 1644511149
transform 1 0 44252 0 1 106624
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_192_475
timestamp 1644511149
transform 1 0 44804 0 1 106624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_192_477
timestamp 1644511149
transform 1 0 44988 0 1 106624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_192_489
timestamp 1644511149
transform 1 0 46092 0 1 106624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_192_501
timestamp 1644511149
transform 1 0 47196 0 1 106624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_192_513
timestamp 1644511149
transform 1 0 48300 0 1 106624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_192_525
timestamp 1644511149
transform 1 0 49404 0 1 106624
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_192_531
timestamp 1644511149
transform 1 0 49956 0 1 106624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_192_533
timestamp 1644511149
transform 1 0 50140 0 1 106624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_192_545
timestamp 1644511149
transform 1 0 51244 0 1 106624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_192_557
timestamp 1644511149
transform 1 0 52348 0 1 106624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_192_569
timestamp 1644511149
transform 1 0 53452 0 1 106624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_192_581
timestamp 1644511149
transform 1 0 54556 0 1 106624
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_192_587
timestamp 1644511149
transform 1 0 55108 0 1 106624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_192_589
timestamp 1644511149
transform 1 0 55292 0 1 106624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_192_601
timestamp 1644511149
transform 1 0 56396 0 1 106624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_192_613
timestamp 1644511149
transform 1 0 57500 0 1 106624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_192_625
timestamp 1644511149
transform 1 0 58604 0 1 106624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_192_637
timestamp 1644511149
transform 1 0 59708 0 1 106624
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_192_643
timestamp 1644511149
transform 1 0 60260 0 1 106624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_192_645
timestamp 1644511149
transform 1 0 60444 0 1 106624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_192_657
timestamp 1644511149
transform 1 0 61548 0 1 106624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_192_669
timestamp 1644511149
transform 1 0 62652 0 1 106624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_192_681
timestamp 1644511149
transform 1 0 63756 0 1 106624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_192_693
timestamp 1644511149
transform 1 0 64860 0 1 106624
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_192_699
timestamp 1644511149
transform 1 0 65412 0 1 106624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_192_701
timestamp 1644511149
transform 1 0 65596 0 1 106624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_192_713
timestamp 1644511149
transform 1 0 66700 0 1 106624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_192_725
timestamp 1644511149
transform 1 0 67804 0 1 106624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_192_737
timestamp 1644511149
transform 1 0 68908 0 1 106624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_192_749
timestamp 1644511149
transform 1 0 70012 0 1 106624
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_192_755
timestamp 1644511149
transform 1 0 70564 0 1 106624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_192_757
timestamp 1644511149
transform 1 0 70748 0 1 106624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_192_769
timestamp 1644511149
transform 1 0 71852 0 1 106624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_192_781
timestamp 1644511149
transform 1 0 72956 0 1 106624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_192_793
timestamp 1644511149
transform 1 0 74060 0 1 106624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_192_805
timestamp 1644511149
transform 1 0 75164 0 1 106624
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_192_811
timestamp 1644511149
transform 1 0 75716 0 1 106624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_192_813
timestamp 1644511149
transform 1 0 75900 0 1 106624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_192_825
timestamp 1644511149
transform 1 0 77004 0 1 106624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_192_837
timestamp 1644511149
transform 1 0 78108 0 1 106624
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_192_841
timestamp 1644511149
transform 1 0 78476 0 1 106624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_193_3
timestamp 1644511149
transform 1 0 1380 0 -1 107712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_193_15
timestamp 1644511149
transform 1 0 2484 0 -1 107712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_193_27
timestamp 1644511149
transform 1 0 3588 0 -1 107712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_193_39
timestamp 1644511149
transform 1 0 4692 0 -1 107712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_193_51
timestamp 1644511149
transform 1 0 5796 0 -1 107712
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_193_55
timestamp 1644511149
transform 1 0 6164 0 -1 107712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_193_57
timestamp 1644511149
transform 1 0 6348 0 -1 107712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_193_69
timestamp 1644511149
transform 1 0 7452 0 -1 107712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_193_81
timestamp 1644511149
transform 1 0 8556 0 -1 107712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_193_93
timestamp 1644511149
transform 1 0 9660 0 -1 107712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_193_105
timestamp 1644511149
transform 1 0 10764 0 -1 107712
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_193_111
timestamp 1644511149
transform 1 0 11316 0 -1 107712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_193_113
timestamp 1644511149
transform 1 0 11500 0 -1 107712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_193_125
timestamp 1644511149
transform 1 0 12604 0 -1 107712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_193_137
timestamp 1644511149
transform 1 0 13708 0 -1 107712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_193_149
timestamp 1644511149
transform 1 0 14812 0 -1 107712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_193_161
timestamp 1644511149
transform 1 0 15916 0 -1 107712
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_193_167
timestamp 1644511149
transform 1 0 16468 0 -1 107712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_193_169
timestamp 1644511149
transform 1 0 16652 0 -1 107712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_193_181
timestamp 1644511149
transform 1 0 17756 0 -1 107712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_193_193
timestamp 1644511149
transform 1 0 18860 0 -1 107712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_193_205
timestamp 1644511149
transform 1 0 19964 0 -1 107712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_193_217
timestamp 1644511149
transform 1 0 21068 0 -1 107712
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_193_223
timestamp 1644511149
transform 1 0 21620 0 -1 107712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_193_225
timestamp 1644511149
transform 1 0 21804 0 -1 107712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_193_237
timestamp 1644511149
transform 1 0 22908 0 -1 107712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_193_249
timestamp 1644511149
transform 1 0 24012 0 -1 107712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_193_261
timestamp 1644511149
transform 1 0 25116 0 -1 107712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_193_273
timestamp 1644511149
transform 1 0 26220 0 -1 107712
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_193_279
timestamp 1644511149
transform 1 0 26772 0 -1 107712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_193_281
timestamp 1644511149
transform 1 0 26956 0 -1 107712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_193_293
timestamp 1644511149
transform 1 0 28060 0 -1 107712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_193_305
timestamp 1644511149
transform 1 0 29164 0 -1 107712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_193_317
timestamp 1644511149
transform 1 0 30268 0 -1 107712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_193_329
timestamp 1644511149
transform 1 0 31372 0 -1 107712
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_193_335
timestamp 1644511149
transform 1 0 31924 0 -1 107712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_193_337
timestamp 1644511149
transform 1 0 32108 0 -1 107712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_193_349
timestamp 1644511149
transform 1 0 33212 0 -1 107712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_193_361
timestamp 1644511149
transform 1 0 34316 0 -1 107712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_193_373
timestamp 1644511149
transform 1 0 35420 0 -1 107712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_193_385
timestamp 1644511149
transform 1 0 36524 0 -1 107712
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_193_391
timestamp 1644511149
transform 1 0 37076 0 -1 107712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_193_393
timestamp 1644511149
transform 1 0 37260 0 -1 107712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_193_405
timestamp 1644511149
transform 1 0 38364 0 -1 107712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_193_417
timestamp 1644511149
transform 1 0 39468 0 -1 107712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_193_429
timestamp 1644511149
transform 1 0 40572 0 -1 107712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_193_441
timestamp 1644511149
transform 1 0 41676 0 -1 107712
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_193_447
timestamp 1644511149
transform 1 0 42228 0 -1 107712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_193_449
timestamp 1644511149
transform 1 0 42412 0 -1 107712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_193_461
timestamp 1644511149
transform 1 0 43516 0 -1 107712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_193_473
timestamp 1644511149
transform 1 0 44620 0 -1 107712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_193_485
timestamp 1644511149
transform 1 0 45724 0 -1 107712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_193_497
timestamp 1644511149
transform 1 0 46828 0 -1 107712
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_193_503
timestamp 1644511149
transform 1 0 47380 0 -1 107712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_193_505
timestamp 1644511149
transform 1 0 47564 0 -1 107712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_193_517
timestamp 1644511149
transform 1 0 48668 0 -1 107712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_193_529
timestamp 1644511149
transform 1 0 49772 0 -1 107712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_193_541
timestamp 1644511149
transform 1 0 50876 0 -1 107712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_193_553
timestamp 1644511149
transform 1 0 51980 0 -1 107712
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_193_559
timestamp 1644511149
transform 1 0 52532 0 -1 107712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_193_561
timestamp 1644511149
transform 1 0 52716 0 -1 107712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_193_573
timestamp 1644511149
transform 1 0 53820 0 -1 107712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_193_585
timestamp 1644511149
transform 1 0 54924 0 -1 107712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_193_597
timestamp 1644511149
transform 1 0 56028 0 -1 107712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_193_609
timestamp 1644511149
transform 1 0 57132 0 -1 107712
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_193_615
timestamp 1644511149
transform 1 0 57684 0 -1 107712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_193_617
timestamp 1644511149
transform 1 0 57868 0 -1 107712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_193_629
timestamp 1644511149
transform 1 0 58972 0 -1 107712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_193_641
timestamp 1644511149
transform 1 0 60076 0 -1 107712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_193_653
timestamp 1644511149
transform 1 0 61180 0 -1 107712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_193_665
timestamp 1644511149
transform 1 0 62284 0 -1 107712
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_193_671
timestamp 1644511149
transform 1 0 62836 0 -1 107712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_193_673
timestamp 1644511149
transform 1 0 63020 0 -1 107712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_193_685
timestamp 1644511149
transform 1 0 64124 0 -1 107712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_193_697
timestamp 1644511149
transform 1 0 65228 0 -1 107712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_193_709
timestamp 1644511149
transform 1 0 66332 0 -1 107712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_193_721
timestamp 1644511149
transform 1 0 67436 0 -1 107712
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_193_727
timestamp 1644511149
transform 1 0 67988 0 -1 107712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_193_729
timestamp 1644511149
transform 1 0 68172 0 -1 107712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_193_741
timestamp 1644511149
transform 1 0 69276 0 -1 107712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_193_753
timestamp 1644511149
transform 1 0 70380 0 -1 107712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_193_765
timestamp 1644511149
transform 1 0 71484 0 -1 107712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_193_777
timestamp 1644511149
transform 1 0 72588 0 -1 107712
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_193_783
timestamp 1644511149
transform 1 0 73140 0 -1 107712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_193_785
timestamp 1644511149
transform 1 0 73324 0 -1 107712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_193_797
timestamp 1644511149
transform 1 0 74428 0 -1 107712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_193_809
timestamp 1644511149
transform 1 0 75532 0 -1 107712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_193_821
timestamp 1644511149
transform 1 0 76636 0 -1 107712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_193_833
timestamp 1644511149
transform 1 0 77740 0 -1 107712
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_193_839
timestamp 1644511149
transform 1 0 78292 0 -1 107712
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_193_841
timestamp 1644511149
transform 1 0 78476 0 -1 107712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_194_3
timestamp 1644511149
transform 1 0 1380 0 1 107712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_194_15
timestamp 1644511149
transform 1 0 2484 0 1 107712
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_194_27
timestamp 1644511149
transform 1 0 3588 0 1 107712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_194_29
timestamp 1644511149
transform 1 0 3772 0 1 107712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_194_41
timestamp 1644511149
transform 1 0 4876 0 1 107712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_194_53
timestamp 1644511149
transform 1 0 5980 0 1 107712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_194_65
timestamp 1644511149
transform 1 0 7084 0 1 107712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_194_77
timestamp 1644511149
transform 1 0 8188 0 1 107712
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_194_83
timestamp 1644511149
transform 1 0 8740 0 1 107712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_194_85
timestamp 1644511149
transform 1 0 8924 0 1 107712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_194_97
timestamp 1644511149
transform 1 0 10028 0 1 107712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_194_109
timestamp 1644511149
transform 1 0 11132 0 1 107712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_194_121
timestamp 1644511149
transform 1 0 12236 0 1 107712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_194_133
timestamp 1644511149
transform 1 0 13340 0 1 107712
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_194_139
timestamp 1644511149
transform 1 0 13892 0 1 107712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_194_141
timestamp 1644511149
transform 1 0 14076 0 1 107712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_194_153
timestamp 1644511149
transform 1 0 15180 0 1 107712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_194_165
timestamp 1644511149
transform 1 0 16284 0 1 107712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_194_177
timestamp 1644511149
transform 1 0 17388 0 1 107712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_194_189
timestamp 1644511149
transform 1 0 18492 0 1 107712
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_194_195
timestamp 1644511149
transform 1 0 19044 0 1 107712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_194_197
timestamp 1644511149
transform 1 0 19228 0 1 107712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_194_209
timestamp 1644511149
transform 1 0 20332 0 1 107712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_194_221
timestamp 1644511149
transform 1 0 21436 0 1 107712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_194_233
timestamp 1644511149
transform 1 0 22540 0 1 107712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_194_245
timestamp 1644511149
transform 1 0 23644 0 1 107712
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_194_251
timestamp 1644511149
transform 1 0 24196 0 1 107712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_194_253
timestamp 1644511149
transform 1 0 24380 0 1 107712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_194_265
timestamp 1644511149
transform 1 0 25484 0 1 107712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_194_277
timestamp 1644511149
transform 1 0 26588 0 1 107712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_194_289
timestamp 1644511149
transform 1 0 27692 0 1 107712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_194_301
timestamp 1644511149
transform 1 0 28796 0 1 107712
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_194_307
timestamp 1644511149
transform 1 0 29348 0 1 107712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_194_309
timestamp 1644511149
transform 1 0 29532 0 1 107712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_194_321
timestamp 1644511149
transform 1 0 30636 0 1 107712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_194_333
timestamp 1644511149
transform 1 0 31740 0 1 107712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_194_345
timestamp 1644511149
transform 1 0 32844 0 1 107712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_194_357
timestamp 1644511149
transform 1 0 33948 0 1 107712
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_194_363
timestamp 1644511149
transform 1 0 34500 0 1 107712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_194_365
timestamp 1644511149
transform 1 0 34684 0 1 107712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_194_377
timestamp 1644511149
transform 1 0 35788 0 1 107712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_194_389
timestamp 1644511149
transform 1 0 36892 0 1 107712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_194_401
timestamp 1644511149
transform 1 0 37996 0 1 107712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_194_413
timestamp 1644511149
transform 1 0 39100 0 1 107712
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_194_419
timestamp 1644511149
transform 1 0 39652 0 1 107712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_194_421
timestamp 1644511149
transform 1 0 39836 0 1 107712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_194_433
timestamp 1644511149
transform 1 0 40940 0 1 107712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_194_445
timestamp 1644511149
transform 1 0 42044 0 1 107712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_194_457
timestamp 1644511149
transform 1 0 43148 0 1 107712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_194_469
timestamp 1644511149
transform 1 0 44252 0 1 107712
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_194_475
timestamp 1644511149
transform 1 0 44804 0 1 107712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_194_477
timestamp 1644511149
transform 1 0 44988 0 1 107712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_194_489
timestamp 1644511149
transform 1 0 46092 0 1 107712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_194_501
timestamp 1644511149
transform 1 0 47196 0 1 107712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_194_513
timestamp 1644511149
transform 1 0 48300 0 1 107712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_194_525
timestamp 1644511149
transform 1 0 49404 0 1 107712
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_194_531
timestamp 1644511149
transform 1 0 49956 0 1 107712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_194_533
timestamp 1644511149
transform 1 0 50140 0 1 107712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_194_545
timestamp 1644511149
transform 1 0 51244 0 1 107712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_194_557
timestamp 1644511149
transform 1 0 52348 0 1 107712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_194_569
timestamp 1644511149
transform 1 0 53452 0 1 107712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_194_581
timestamp 1644511149
transform 1 0 54556 0 1 107712
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_194_587
timestamp 1644511149
transform 1 0 55108 0 1 107712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_194_589
timestamp 1644511149
transform 1 0 55292 0 1 107712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_194_601
timestamp 1644511149
transform 1 0 56396 0 1 107712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_194_613
timestamp 1644511149
transform 1 0 57500 0 1 107712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_194_625
timestamp 1644511149
transform 1 0 58604 0 1 107712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_194_637
timestamp 1644511149
transform 1 0 59708 0 1 107712
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_194_643
timestamp 1644511149
transform 1 0 60260 0 1 107712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_194_645
timestamp 1644511149
transform 1 0 60444 0 1 107712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_194_657
timestamp 1644511149
transform 1 0 61548 0 1 107712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_194_669
timestamp 1644511149
transform 1 0 62652 0 1 107712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_194_681
timestamp 1644511149
transform 1 0 63756 0 1 107712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_194_693
timestamp 1644511149
transform 1 0 64860 0 1 107712
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_194_699
timestamp 1644511149
transform 1 0 65412 0 1 107712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_194_701
timestamp 1644511149
transform 1 0 65596 0 1 107712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_194_713
timestamp 1644511149
transform 1 0 66700 0 1 107712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_194_725
timestamp 1644511149
transform 1 0 67804 0 1 107712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_194_737
timestamp 1644511149
transform 1 0 68908 0 1 107712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_194_749
timestamp 1644511149
transform 1 0 70012 0 1 107712
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_194_755
timestamp 1644511149
transform 1 0 70564 0 1 107712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_194_757
timestamp 1644511149
transform 1 0 70748 0 1 107712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_194_769
timestamp 1644511149
transform 1 0 71852 0 1 107712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_194_781
timestamp 1644511149
transform 1 0 72956 0 1 107712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_194_793
timestamp 1644511149
transform 1 0 74060 0 1 107712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_194_805
timestamp 1644511149
transform 1 0 75164 0 1 107712
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_194_811
timestamp 1644511149
transform 1 0 75716 0 1 107712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_194_813
timestamp 1644511149
transform 1 0 75900 0 1 107712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_194_825
timestamp 1644511149
transform 1 0 77004 0 1 107712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_194_837
timestamp 1644511149
transform 1 0 78108 0 1 107712
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_194_841
timestamp 1644511149
transform 1 0 78476 0 1 107712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_195_3
timestamp 1644511149
transform 1 0 1380 0 -1 108800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_195_15
timestamp 1644511149
transform 1 0 2484 0 -1 108800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_195_27
timestamp 1644511149
transform 1 0 3588 0 -1 108800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_195_39
timestamp 1644511149
transform 1 0 4692 0 -1 108800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_195_51
timestamp 1644511149
transform 1 0 5796 0 -1 108800
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_195_55
timestamp 1644511149
transform 1 0 6164 0 -1 108800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_195_57
timestamp 1644511149
transform 1 0 6348 0 -1 108800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_195_69
timestamp 1644511149
transform 1 0 7452 0 -1 108800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_195_81
timestamp 1644511149
transform 1 0 8556 0 -1 108800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_195_93
timestamp 1644511149
transform 1 0 9660 0 -1 108800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_195_105
timestamp 1644511149
transform 1 0 10764 0 -1 108800
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_195_111
timestamp 1644511149
transform 1 0 11316 0 -1 108800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_195_113
timestamp 1644511149
transform 1 0 11500 0 -1 108800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_195_125
timestamp 1644511149
transform 1 0 12604 0 -1 108800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_195_137
timestamp 1644511149
transform 1 0 13708 0 -1 108800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_195_149
timestamp 1644511149
transform 1 0 14812 0 -1 108800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_195_161
timestamp 1644511149
transform 1 0 15916 0 -1 108800
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_195_167
timestamp 1644511149
transform 1 0 16468 0 -1 108800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_195_169
timestamp 1644511149
transform 1 0 16652 0 -1 108800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_195_181
timestamp 1644511149
transform 1 0 17756 0 -1 108800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_195_193
timestamp 1644511149
transform 1 0 18860 0 -1 108800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_195_205
timestamp 1644511149
transform 1 0 19964 0 -1 108800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_195_217
timestamp 1644511149
transform 1 0 21068 0 -1 108800
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_195_223
timestamp 1644511149
transform 1 0 21620 0 -1 108800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_195_225
timestamp 1644511149
transform 1 0 21804 0 -1 108800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_195_237
timestamp 1644511149
transform 1 0 22908 0 -1 108800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_195_249
timestamp 1644511149
transform 1 0 24012 0 -1 108800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_195_261
timestamp 1644511149
transform 1 0 25116 0 -1 108800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_195_273
timestamp 1644511149
transform 1 0 26220 0 -1 108800
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_195_279
timestamp 1644511149
transform 1 0 26772 0 -1 108800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_195_281
timestamp 1644511149
transform 1 0 26956 0 -1 108800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_195_293
timestamp 1644511149
transform 1 0 28060 0 -1 108800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_195_305
timestamp 1644511149
transform 1 0 29164 0 -1 108800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_195_317
timestamp 1644511149
transform 1 0 30268 0 -1 108800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_195_329
timestamp 1644511149
transform 1 0 31372 0 -1 108800
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_195_335
timestamp 1644511149
transform 1 0 31924 0 -1 108800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_195_337
timestamp 1644511149
transform 1 0 32108 0 -1 108800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_195_349
timestamp 1644511149
transform 1 0 33212 0 -1 108800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_195_361
timestamp 1644511149
transform 1 0 34316 0 -1 108800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_195_373
timestamp 1644511149
transform 1 0 35420 0 -1 108800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_195_385
timestamp 1644511149
transform 1 0 36524 0 -1 108800
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_195_391
timestamp 1644511149
transform 1 0 37076 0 -1 108800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_195_393
timestamp 1644511149
transform 1 0 37260 0 -1 108800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_195_405
timestamp 1644511149
transform 1 0 38364 0 -1 108800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_195_417
timestamp 1644511149
transform 1 0 39468 0 -1 108800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_195_429
timestamp 1644511149
transform 1 0 40572 0 -1 108800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_195_441
timestamp 1644511149
transform 1 0 41676 0 -1 108800
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_195_447
timestamp 1644511149
transform 1 0 42228 0 -1 108800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_195_449
timestamp 1644511149
transform 1 0 42412 0 -1 108800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_195_461
timestamp 1644511149
transform 1 0 43516 0 -1 108800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_195_473
timestamp 1644511149
transform 1 0 44620 0 -1 108800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_195_485
timestamp 1644511149
transform 1 0 45724 0 -1 108800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_195_497
timestamp 1644511149
transform 1 0 46828 0 -1 108800
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_195_503
timestamp 1644511149
transform 1 0 47380 0 -1 108800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_195_505
timestamp 1644511149
transform 1 0 47564 0 -1 108800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_195_517
timestamp 1644511149
transform 1 0 48668 0 -1 108800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_195_529
timestamp 1644511149
transform 1 0 49772 0 -1 108800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_195_541
timestamp 1644511149
transform 1 0 50876 0 -1 108800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_195_553
timestamp 1644511149
transform 1 0 51980 0 -1 108800
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_195_559
timestamp 1644511149
transform 1 0 52532 0 -1 108800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_195_561
timestamp 1644511149
transform 1 0 52716 0 -1 108800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_195_573
timestamp 1644511149
transform 1 0 53820 0 -1 108800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_195_585
timestamp 1644511149
transform 1 0 54924 0 -1 108800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_195_597
timestamp 1644511149
transform 1 0 56028 0 -1 108800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_195_609
timestamp 1644511149
transform 1 0 57132 0 -1 108800
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_195_615
timestamp 1644511149
transform 1 0 57684 0 -1 108800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_195_617
timestamp 1644511149
transform 1 0 57868 0 -1 108800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_195_629
timestamp 1644511149
transform 1 0 58972 0 -1 108800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_195_641
timestamp 1644511149
transform 1 0 60076 0 -1 108800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_195_653
timestamp 1644511149
transform 1 0 61180 0 -1 108800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_195_665
timestamp 1644511149
transform 1 0 62284 0 -1 108800
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_195_671
timestamp 1644511149
transform 1 0 62836 0 -1 108800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_195_673
timestamp 1644511149
transform 1 0 63020 0 -1 108800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_195_685
timestamp 1644511149
transform 1 0 64124 0 -1 108800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_195_697
timestamp 1644511149
transform 1 0 65228 0 -1 108800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_195_709
timestamp 1644511149
transform 1 0 66332 0 -1 108800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_195_721
timestamp 1644511149
transform 1 0 67436 0 -1 108800
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_195_727
timestamp 1644511149
transform 1 0 67988 0 -1 108800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_195_729
timestamp 1644511149
transform 1 0 68172 0 -1 108800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_195_741
timestamp 1644511149
transform 1 0 69276 0 -1 108800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_195_753
timestamp 1644511149
transform 1 0 70380 0 -1 108800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_195_765
timestamp 1644511149
transform 1 0 71484 0 -1 108800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_195_777
timestamp 1644511149
transform 1 0 72588 0 -1 108800
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_195_783
timestamp 1644511149
transform 1 0 73140 0 -1 108800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_195_785
timestamp 1644511149
transform 1 0 73324 0 -1 108800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_195_797
timestamp 1644511149
transform 1 0 74428 0 -1 108800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_195_809
timestamp 1644511149
transform 1 0 75532 0 -1 108800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_195_821
timestamp 1644511149
transform 1 0 76636 0 -1 108800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_195_833
timestamp 1644511149
transform 1 0 77740 0 -1 108800
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_195_839
timestamp 1644511149
transform 1 0 78292 0 -1 108800
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_195_841
timestamp 1644511149
transform 1 0 78476 0 -1 108800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_196_3
timestamp 1644511149
transform 1 0 1380 0 1 108800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_196_15
timestamp 1644511149
transform 1 0 2484 0 1 108800
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_196_27
timestamp 1644511149
transform 1 0 3588 0 1 108800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_196_29
timestamp 1644511149
transform 1 0 3772 0 1 108800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_196_41
timestamp 1644511149
transform 1 0 4876 0 1 108800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_196_53
timestamp 1644511149
transform 1 0 5980 0 1 108800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_196_65
timestamp 1644511149
transform 1 0 7084 0 1 108800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_196_77
timestamp 1644511149
transform 1 0 8188 0 1 108800
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_196_83
timestamp 1644511149
transform 1 0 8740 0 1 108800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_196_85
timestamp 1644511149
transform 1 0 8924 0 1 108800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_196_97
timestamp 1644511149
transform 1 0 10028 0 1 108800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_196_109
timestamp 1644511149
transform 1 0 11132 0 1 108800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_196_121
timestamp 1644511149
transform 1 0 12236 0 1 108800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_196_133
timestamp 1644511149
transform 1 0 13340 0 1 108800
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_196_139
timestamp 1644511149
transform 1 0 13892 0 1 108800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_196_141
timestamp 1644511149
transform 1 0 14076 0 1 108800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_196_153
timestamp 1644511149
transform 1 0 15180 0 1 108800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_196_165
timestamp 1644511149
transform 1 0 16284 0 1 108800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_196_177
timestamp 1644511149
transform 1 0 17388 0 1 108800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_196_189
timestamp 1644511149
transform 1 0 18492 0 1 108800
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_196_195
timestamp 1644511149
transform 1 0 19044 0 1 108800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_196_197
timestamp 1644511149
transform 1 0 19228 0 1 108800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_196_209
timestamp 1644511149
transform 1 0 20332 0 1 108800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_196_221
timestamp 1644511149
transform 1 0 21436 0 1 108800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_196_233
timestamp 1644511149
transform 1 0 22540 0 1 108800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_196_245
timestamp 1644511149
transform 1 0 23644 0 1 108800
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_196_251
timestamp 1644511149
transform 1 0 24196 0 1 108800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_196_253
timestamp 1644511149
transform 1 0 24380 0 1 108800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_196_265
timestamp 1644511149
transform 1 0 25484 0 1 108800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_196_277
timestamp 1644511149
transform 1 0 26588 0 1 108800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_196_289
timestamp 1644511149
transform 1 0 27692 0 1 108800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_196_301
timestamp 1644511149
transform 1 0 28796 0 1 108800
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_196_307
timestamp 1644511149
transform 1 0 29348 0 1 108800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_196_309
timestamp 1644511149
transform 1 0 29532 0 1 108800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_196_321
timestamp 1644511149
transform 1 0 30636 0 1 108800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_196_333
timestamp 1644511149
transform 1 0 31740 0 1 108800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_196_345
timestamp 1644511149
transform 1 0 32844 0 1 108800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_196_357
timestamp 1644511149
transform 1 0 33948 0 1 108800
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_196_363
timestamp 1644511149
transform 1 0 34500 0 1 108800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_196_365
timestamp 1644511149
transform 1 0 34684 0 1 108800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_196_377
timestamp 1644511149
transform 1 0 35788 0 1 108800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_196_389
timestamp 1644511149
transform 1 0 36892 0 1 108800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_196_401
timestamp 1644511149
transform 1 0 37996 0 1 108800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_196_413
timestamp 1644511149
transform 1 0 39100 0 1 108800
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_196_419
timestamp 1644511149
transform 1 0 39652 0 1 108800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_196_425
timestamp 1644511149
transform 1 0 40204 0 1 108800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_196_437
timestamp 1644511149
transform 1 0 41308 0 1 108800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_196_449
timestamp 1644511149
transform 1 0 42412 0 1 108800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_196_461
timestamp 1644511149
transform 1 0 43516 0 1 108800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_196_473
timestamp 1644511149
transform 1 0 44620 0 1 108800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_196_477
timestamp 1644511149
transform 1 0 44988 0 1 108800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_196_489
timestamp 1644511149
transform 1 0 46092 0 1 108800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_196_501
timestamp 1644511149
transform 1 0 47196 0 1 108800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_196_513
timestamp 1644511149
transform 1 0 48300 0 1 108800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_196_525
timestamp 1644511149
transform 1 0 49404 0 1 108800
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_196_531
timestamp 1644511149
transform 1 0 49956 0 1 108800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_196_533
timestamp 1644511149
transform 1 0 50140 0 1 108800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_196_545
timestamp 1644511149
transform 1 0 51244 0 1 108800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_196_557
timestamp 1644511149
transform 1 0 52348 0 1 108800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_196_569
timestamp 1644511149
transform 1 0 53452 0 1 108800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_196_581
timestamp 1644511149
transform 1 0 54556 0 1 108800
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_196_587
timestamp 1644511149
transform 1 0 55108 0 1 108800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_196_589
timestamp 1644511149
transform 1 0 55292 0 1 108800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_196_601
timestamp 1644511149
transform 1 0 56396 0 1 108800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_196_613
timestamp 1644511149
transform 1 0 57500 0 1 108800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_196_625
timestamp 1644511149
transform 1 0 58604 0 1 108800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_196_637
timestamp 1644511149
transform 1 0 59708 0 1 108800
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_196_643
timestamp 1644511149
transform 1 0 60260 0 1 108800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_196_645
timestamp 1644511149
transform 1 0 60444 0 1 108800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_196_657
timestamp 1644511149
transform 1 0 61548 0 1 108800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_196_669
timestamp 1644511149
transform 1 0 62652 0 1 108800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_196_681
timestamp 1644511149
transform 1 0 63756 0 1 108800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_196_693
timestamp 1644511149
transform 1 0 64860 0 1 108800
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_196_699
timestamp 1644511149
transform 1 0 65412 0 1 108800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_196_701
timestamp 1644511149
transform 1 0 65596 0 1 108800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_196_713
timestamp 1644511149
transform 1 0 66700 0 1 108800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_196_725
timestamp 1644511149
transform 1 0 67804 0 1 108800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_196_737
timestamp 1644511149
transform 1 0 68908 0 1 108800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_196_749
timestamp 1644511149
transform 1 0 70012 0 1 108800
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_196_755
timestamp 1644511149
transform 1 0 70564 0 1 108800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_196_757
timestamp 1644511149
transform 1 0 70748 0 1 108800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_196_769
timestamp 1644511149
transform 1 0 71852 0 1 108800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_196_781
timestamp 1644511149
transform 1 0 72956 0 1 108800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_196_793
timestamp 1644511149
transform 1 0 74060 0 1 108800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_196_805
timestamp 1644511149
transform 1 0 75164 0 1 108800
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_196_811
timestamp 1644511149
transform 1 0 75716 0 1 108800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_196_813
timestamp 1644511149
transform 1 0 75900 0 1 108800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_196_825
timestamp 1644511149
transform 1 0 77004 0 1 108800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_196_837
timestamp 1644511149
transform 1 0 78108 0 1 108800
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_196_841
timestamp 1644511149
transform 1 0 78476 0 1 108800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_197_3
timestamp 1644511149
transform 1 0 1380 0 -1 109888
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_197_11
timestamp 1644511149
transform 1 0 2116 0 -1 109888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_197_23
timestamp 1644511149
transform 1 0 3220 0 -1 109888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_197_35
timestamp 1644511149
transform 1 0 4324 0 -1 109888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_197_47
timestamp 1644511149
transform 1 0 5428 0 -1 109888
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_197_55
timestamp 1644511149
transform 1 0 6164 0 -1 109888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_197_57
timestamp 1644511149
transform 1 0 6348 0 -1 109888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_197_69
timestamp 1644511149
transform 1 0 7452 0 -1 109888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_197_81
timestamp 1644511149
transform 1 0 8556 0 -1 109888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_197_93
timestamp 1644511149
transform 1 0 9660 0 -1 109888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_197_105
timestamp 1644511149
transform 1 0 10764 0 -1 109888
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_197_111
timestamp 1644511149
transform 1 0 11316 0 -1 109888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_197_113
timestamp 1644511149
transform 1 0 11500 0 -1 109888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_197_125
timestamp 1644511149
transform 1 0 12604 0 -1 109888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_197_137
timestamp 1644511149
transform 1 0 13708 0 -1 109888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_197_149
timestamp 1644511149
transform 1 0 14812 0 -1 109888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_197_161
timestamp 1644511149
transform 1 0 15916 0 -1 109888
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_197_167
timestamp 1644511149
transform 1 0 16468 0 -1 109888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_197_169
timestamp 1644511149
transform 1 0 16652 0 -1 109888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_197_181
timestamp 1644511149
transform 1 0 17756 0 -1 109888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_197_193
timestamp 1644511149
transform 1 0 18860 0 -1 109888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_197_205
timestamp 1644511149
transform 1 0 19964 0 -1 109888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_197_217
timestamp 1644511149
transform 1 0 21068 0 -1 109888
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_197_223
timestamp 1644511149
transform 1 0 21620 0 -1 109888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_197_225
timestamp 1644511149
transform 1 0 21804 0 -1 109888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_197_237
timestamp 1644511149
transform 1 0 22908 0 -1 109888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_197_249
timestamp 1644511149
transform 1 0 24012 0 -1 109888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_197_261
timestamp 1644511149
transform 1 0 25116 0 -1 109888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_197_273
timestamp 1644511149
transform 1 0 26220 0 -1 109888
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_197_279
timestamp 1644511149
transform 1 0 26772 0 -1 109888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_197_281
timestamp 1644511149
transform 1 0 26956 0 -1 109888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_197_293
timestamp 1644511149
transform 1 0 28060 0 -1 109888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_197_305
timestamp 1644511149
transform 1 0 29164 0 -1 109888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_197_317
timestamp 1644511149
transform 1 0 30268 0 -1 109888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_197_329
timestamp 1644511149
transform 1 0 31372 0 -1 109888
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_197_335
timestamp 1644511149
transform 1 0 31924 0 -1 109888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_197_337
timestamp 1644511149
transform 1 0 32108 0 -1 109888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_197_349
timestamp 1644511149
transform 1 0 33212 0 -1 109888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_197_361
timestamp 1644511149
transform 1 0 34316 0 -1 109888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_197_373
timestamp 1644511149
transform 1 0 35420 0 -1 109888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_197_385
timestamp 1644511149
transform 1 0 36524 0 -1 109888
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_197_391
timestamp 1644511149
transform 1 0 37076 0 -1 109888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_197_393
timestamp 1644511149
transform 1 0 37260 0 -1 109888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_197_405
timestamp 1644511149
transform 1 0 38364 0 -1 109888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_197_417
timestamp 1644511149
transform 1 0 39468 0 -1 109888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_197_429
timestamp 1644511149
transform 1 0 40572 0 -1 109888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_197_441
timestamp 1644511149
transform 1 0 41676 0 -1 109888
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_197_447
timestamp 1644511149
transform 1 0 42228 0 -1 109888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_197_449
timestamp 1644511149
transform 1 0 42412 0 -1 109888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_197_461
timestamp 1644511149
transform 1 0 43516 0 -1 109888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_197_473
timestamp 1644511149
transform 1 0 44620 0 -1 109888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_197_485
timestamp 1644511149
transform 1 0 45724 0 -1 109888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_197_497
timestamp 1644511149
transform 1 0 46828 0 -1 109888
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_197_503
timestamp 1644511149
transform 1 0 47380 0 -1 109888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_197_505
timestamp 1644511149
transform 1 0 47564 0 -1 109888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_197_517
timestamp 1644511149
transform 1 0 48668 0 -1 109888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_197_529
timestamp 1644511149
transform 1 0 49772 0 -1 109888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_197_541
timestamp 1644511149
transform 1 0 50876 0 -1 109888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_197_553
timestamp 1644511149
transform 1 0 51980 0 -1 109888
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_197_559
timestamp 1644511149
transform 1 0 52532 0 -1 109888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_197_561
timestamp 1644511149
transform 1 0 52716 0 -1 109888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_197_573
timestamp 1644511149
transform 1 0 53820 0 -1 109888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_197_585
timestamp 1644511149
transform 1 0 54924 0 -1 109888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_197_597
timestamp 1644511149
transform 1 0 56028 0 -1 109888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_197_609
timestamp 1644511149
transform 1 0 57132 0 -1 109888
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_197_615
timestamp 1644511149
transform 1 0 57684 0 -1 109888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_197_617
timestamp 1644511149
transform 1 0 57868 0 -1 109888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_197_629
timestamp 1644511149
transform 1 0 58972 0 -1 109888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_197_641
timestamp 1644511149
transform 1 0 60076 0 -1 109888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_197_653
timestamp 1644511149
transform 1 0 61180 0 -1 109888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_197_665
timestamp 1644511149
transform 1 0 62284 0 -1 109888
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_197_671
timestamp 1644511149
transform 1 0 62836 0 -1 109888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_197_673
timestamp 1644511149
transform 1 0 63020 0 -1 109888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_197_685
timestamp 1644511149
transform 1 0 64124 0 -1 109888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_197_697
timestamp 1644511149
transform 1 0 65228 0 -1 109888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_197_709
timestamp 1644511149
transform 1 0 66332 0 -1 109888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_197_721
timestamp 1644511149
transform 1 0 67436 0 -1 109888
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_197_727
timestamp 1644511149
transform 1 0 67988 0 -1 109888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_197_729
timestamp 1644511149
transform 1 0 68172 0 -1 109888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_197_741
timestamp 1644511149
transform 1 0 69276 0 -1 109888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_197_753
timestamp 1644511149
transform 1 0 70380 0 -1 109888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_197_765
timestamp 1644511149
transform 1 0 71484 0 -1 109888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_197_777
timestamp 1644511149
transform 1 0 72588 0 -1 109888
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_197_783
timestamp 1644511149
transform 1 0 73140 0 -1 109888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_197_785
timestamp 1644511149
transform 1 0 73324 0 -1 109888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_197_797
timestamp 1644511149
transform 1 0 74428 0 -1 109888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_197_809
timestamp 1644511149
transform 1 0 75532 0 -1 109888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_197_821
timestamp 1644511149
transform 1 0 76636 0 -1 109888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_197_833
timestamp 1644511149
transform 1 0 77740 0 -1 109888
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_197_839
timestamp 1644511149
transform 1 0 78292 0 -1 109888
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_197_841
timestamp 1644511149
transform 1 0 78476 0 -1 109888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_198_3
timestamp 1644511149
transform 1 0 1380 0 1 109888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_198_15
timestamp 1644511149
transform 1 0 2484 0 1 109888
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_198_27
timestamp 1644511149
transform 1 0 3588 0 1 109888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_198_29
timestamp 1644511149
transform 1 0 3772 0 1 109888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_198_41
timestamp 1644511149
transform 1 0 4876 0 1 109888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_198_53
timestamp 1644511149
transform 1 0 5980 0 1 109888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_198_65
timestamp 1644511149
transform 1 0 7084 0 1 109888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_198_77
timestamp 1644511149
transform 1 0 8188 0 1 109888
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_198_83
timestamp 1644511149
transform 1 0 8740 0 1 109888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_198_85
timestamp 1644511149
transform 1 0 8924 0 1 109888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_198_97
timestamp 1644511149
transform 1 0 10028 0 1 109888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_198_109
timestamp 1644511149
transform 1 0 11132 0 1 109888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_198_121
timestamp 1644511149
transform 1 0 12236 0 1 109888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_198_133
timestamp 1644511149
transform 1 0 13340 0 1 109888
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_198_139
timestamp 1644511149
transform 1 0 13892 0 1 109888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_198_141
timestamp 1644511149
transform 1 0 14076 0 1 109888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_198_153
timestamp 1644511149
transform 1 0 15180 0 1 109888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_198_165
timestamp 1644511149
transform 1 0 16284 0 1 109888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_198_177
timestamp 1644511149
transform 1 0 17388 0 1 109888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_198_189
timestamp 1644511149
transform 1 0 18492 0 1 109888
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_198_195
timestamp 1644511149
transform 1 0 19044 0 1 109888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_198_197
timestamp 1644511149
transform 1 0 19228 0 1 109888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_198_209
timestamp 1644511149
transform 1 0 20332 0 1 109888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_198_221
timestamp 1644511149
transform 1 0 21436 0 1 109888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_198_233
timestamp 1644511149
transform 1 0 22540 0 1 109888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_198_245
timestamp 1644511149
transform 1 0 23644 0 1 109888
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_198_251
timestamp 1644511149
transform 1 0 24196 0 1 109888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_198_253
timestamp 1644511149
transform 1 0 24380 0 1 109888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_198_265
timestamp 1644511149
transform 1 0 25484 0 1 109888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_198_277
timestamp 1644511149
transform 1 0 26588 0 1 109888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_198_289
timestamp 1644511149
transform 1 0 27692 0 1 109888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_198_301
timestamp 1644511149
transform 1 0 28796 0 1 109888
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_198_307
timestamp 1644511149
transform 1 0 29348 0 1 109888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_198_309
timestamp 1644511149
transform 1 0 29532 0 1 109888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_198_321
timestamp 1644511149
transform 1 0 30636 0 1 109888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_198_333
timestamp 1644511149
transform 1 0 31740 0 1 109888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_198_345
timestamp 1644511149
transform 1 0 32844 0 1 109888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_198_357
timestamp 1644511149
transform 1 0 33948 0 1 109888
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_198_363
timestamp 1644511149
transform 1 0 34500 0 1 109888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_198_365
timestamp 1644511149
transform 1 0 34684 0 1 109888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_198_377
timestamp 1644511149
transform 1 0 35788 0 1 109888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_198_389
timestamp 1644511149
transform 1 0 36892 0 1 109888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_198_401
timestamp 1644511149
transform 1 0 37996 0 1 109888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_198_413
timestamp 1644511149
transform 1 0 39100 0 1 109888
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_198_419
timestamp 1644511149
transform 1 0 39652 0 1 109888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_198_421
timestamp 1644511149
transform 1 0 39836 0 1 109888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_198_433
timestamp 1644511149
transform 1 0 40940 0 1 109888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_198_445
timestamp 1644511149
transform 1 0 42044 0 1 109888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_198_457
timestamp 1644511149
transform 1 0 43148 0 1 109888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_198_469
timestamp 1644511149
transform 1 0 44252 0 1 109888
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_198_475
timestamp 1644511149
transform 1 0 44804 0 1 109888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_198_477
timestamp 1644511149
transform 1 0 44988 0 1 109888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_198_489
timestamp 1644511149
transform 1 0 46092 0 1 109888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_198_501
timestamp 1644511149
transform 1 0 47196 0 1 109888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_198_513
timestamp 1644511149
transform 1 0 48300 0 1 109888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_198_525
timestamp 1644511149
transform 1 0 49404 0 1 109888
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_198_531
timestamp 1644511149
transform 1 0 49956 0 1 109888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_198_533
timestamp 1644511149
transform 1 0 50140 0 1 109888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_198_545
timestamp 1644511149
transform 1 0 51244 0 1 109888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_198_557
timestamp 1644511149
transform 1 0 52348 0 1 109888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_198_569
timestamp 1644511149
transform 1 0 53452 0 1 109888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_198_581
timestamp 1644511149
transform 1 0 54556 0 1 109888
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_198_587
timestamp 1644511149
transform 1 0 55108 0 1 109888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_198_589
timestamp 1644511149
transform 1 0 55292 0 1 109888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_198_601
timestamp 1644511149
transform 1 0 56396 0 1 109888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_198_613
timestamp 1644511149
transform 1 0 57500 0 1 109888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_198_625
timestamp 1644511149
transform 1 0 58604 0 1 109888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_198_637
timestamp 1644511149
transform 1 0 59708 0 1 109888
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_198_643
timestamp 1644511149
transform 1 0 60260 0 1 109888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_198_645
timestamp 1644511149
transform 1 0 60444 0 1 109888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_198_657
timestamp 1644511149
transform 1 0 61548 0 1 109888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_198_669
timestamp 1644511149
transform 1 0 62652 0 1 109888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_198_681
timestamp 1644511149
transform 1 0 63756 0 1 109888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_198_693
timestamp 1644511149
transform 1 0 64860 0 1 109888
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_198_699
timestamp 1644511149
transform 1 0 65412 0 1 109888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_198_701
timestamp 1644511149
transform 1 0 65596 0 1 109888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_198_713
timestamp 1644511149
transform 1 0 66700 0 1 109888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_198_725
timestamp 1644511149
transform 1 0 67804 0 1 109888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_198_737
timestamp 1644511149
transform 1 0 68908 0 1 109888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_198_749
timestamp 1644511149
transform 1 0 70012 0 1 109888
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_198_755
timestamp 1644511149
transform 1 0 70564 0 1 109888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_198_757
timestamp 1644511149
transform 1 0 70748 0 1 109888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_198_769
timestamp 1644511149
transform 1 0 71852 0 1 109888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_198_781
timestamp 1644511149
transform 1 0 72956 0 1 109888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_198_793
timestamp 1644511149
transform 1 0 74060 0 1 109888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_198_805
timestamp 1644511149
transform 1 0 75164 0 1 109888
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_198_811
timestamp 1644511149
transform 1 0 75716 0 1 109888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_198_813
timestamp 1644511149
transform 1 0 75900 0 1 109888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_198_825
timestamp 1644511149
transform 1 0 77004 0 1 109888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_198_837
timestamp 1644511149
transform 1 0 78108 0 1 109888
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_198_841
timestamp 1644511149
transform 1 0 78476 0 1 109888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_199_3
timestamp 1644511149
transform 1 0 1380 0 -1 110976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_199_15
timestamp 1644511149
transform 1 0 2484 0 -1 110976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_199_27
timestamp 1644511149
transform 1 0 3588 0 -1 110976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_199_39
timestamp 1644511149
transform 1 0 4692 0 -1 110976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_199_51
timestamp 1644511149
transform 1 0 5796 0 -1 110976
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_199_55
timestamp 1644511149
transform 1 0 6164 0 -1 110976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_199_57
timestamp 1644511149
transform 1 0 6348 0 -1 110976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_199_69
timestamp 1644511149
transform 1 0 7452 0 -1 110976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_199_81
timestamp 1644511149
transform 1 0 8556 0 -1 110976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_199_93
timestamp 1644511149
transform 1 0 9660 0 -1 110976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_199_105
timestamp 1644511149
transform 1 0 10764 0 -1 110976
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_199_111
timestamp 1644511149
transform 1 0 11316 0 -1 110976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_199_113
timestamp 1644511149
transform 1 0 11500 0 -1 110976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_199_125
timestamp 1644511149
transform 1 0 12604 0 -1 110976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_199_137
timestamp 1644511149
transform 1 0 13708 0 -1 110976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_199_149
timestamp 1644511149
transform 1 0 14812 0 -1 110976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_199_161
timestamp 1644511149
transform 1 0 15916 0 -1 110976
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_199_167
timestamp 1644511149
transform 1 0 16468 0 -1 110976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_199_169
timestamp 1644511149
transform 1 0 16652 0 -1 110976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_199_181
timestamp 1644511149
transform 1 0 17756 0 -1 110976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_199_193
timestamp 1644511149
transform 1 0 18860 0 -1 110976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_199_205
timestamp 1644511149
transform 1 0 19964 0 -1 110976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_199_217
timestamp 1644511149
transform 1 0 21068 0 -1 110976
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_199_223
timestamp 1644511149
transform 1 0 21620 0 -1 110976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_199_225
timestamp 1644511149
transform 1 0 21804 0 -1 110976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_199_237
timestamp 1644511149
transform 1 0 22908 0 -1 110976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_199_249
timestamp 1644511149
transform 1 0 24012 0 -1 110976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_199_261
timestamp 1644511149
transform 1 0 25116 0 -1 110976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_199_273
timestamp 1644511149
transform 1 0 26220 0 -1 110976
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_199_279
timestamp 1644511149
transform 1 0 26772 0 -1 110976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_199_281
timestamp 1644511149
transform 1 0 26956 0 -1 110976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_199_293
timestamp 1644511149
transform 1 0 28060 0 -1 110976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_199_305
timestamp 1644511149
transform 1 0 29164 0 -1 110976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_199_317
timestamp 1644511149
transform 1 0 30268 0 -1 110976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_199_329
timestamp 1644511149
transform 1 0 31372 0 -1 110976
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_199_335
timestamp 1644511149
transform 1 0 31924 0 -1 110976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_199_337
timestamp 1644511149
transform 1 0 32108 0 -1 110976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_199_349
timestamp 1644511149
transform 1 0 33212 0 -1 110976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_199_361
timestamp 1644511149
transform 1 0 34316 0 -1 110976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_199_373
timestamp 1644511149
transform 1 0 35420 0 -1 110976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_199_385
timestamp 1644511149
transform 1 0 36524 0 -1 110976
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_199_391
timestamp 1644511149
transform 1 0 37076 0 -1 110976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_199_393
timestamp 1644511149
transform 1 0 37260 0 -1 110976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_199_405
timestamp 1644511149
transform 1 0 38364 0 -1 110976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_199_417
timestamp 1644511149
transform 1 0 39468 0 -1 110976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_199_429
timestamp 1644511149
transform 1 0 40572 0 -1 110976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_199_441
timestamp 1644511149
transform 1 0 41676 0 -1 110976
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_199_447
timestamp 1644511149
transform 1 0 42228 0 -1 110976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_199_449
timestamp 1644511149
transform 1 0 42412 0 -1 110976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_199_461
timestamp 1644511149
transform 1 0 43516 0 -1 110976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_199_473
timestamp 1644511149
transform 1 0 44620 0 -1 110976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_199_485
timestamp 1644511149
transform 1 0 45724 0 -1 110976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_199_497
timestamp 1644511149
transform 1 0 46828 0 -1 110976
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_199_503
timestamp 1644511149
transform 1 0 47380 0 -1 110976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_199_505
timestamp 1644511149
transform 1 0 47564 0 -1 110976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_199_517
timestamp 1644511149
transform 1 0 48668 0 -1 110976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_199_529
timestamp 1644511149
transform 1 0 49772 0 -1 110976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_199_541
timestamp 1644511149
transform 1 0 50876 0 -1 110976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_199_553
timestamp 1644511149
transform 1 0 51980 0 -1 110976
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_199_559
timestamp 1644511149
transform 1 0 52532 0 -1 110976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_199_561
timestamp 1644511149
transform 1 0 52716 0 -1 110976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_199_573
timestamp 1644511149
transform 1 0 53820 0 -1 110976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_199_585
timestamp 1644511149
transform 1 0 54924 0 -1 110976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_199_597
timestamp 1644511149
transform 1 0 56028 0 -1 110976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_199_609
timestamp 1644511149
transform 1 0 57132 0 -1 110976
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_199_615
timestamp 1644511149
transform 1 0 57684 0 -1 110976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_199_617
timestamp 1644511149
transform 1 0 57868 0 -1 110976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_199_629
timestamp 1644511149
transform 1 0 58972 0 -1 110976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_199_641
timestamp 1644511149
transform 1 0 60076 0 -1 110976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_199_653
timestamp 1644511149
transform 1 0 61180 0 -1 110976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_199_665
timestamp 1644511149
transform 1 0 62284 0 -1 110976
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_199_671
timestamp 1644511149
transform 1 0 62836 0 -1 110976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_199_673
timestamp 1644511149
transform 1 0 63020 0 -1 110976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_199_685
timestamp 1644511149
transform 1 0 64124 0 -1 110976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_199_697
timestamp 1644511149
transform 1 0 65228 0 -1 110976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_199_709
timestamp 1644511149
transform 1 0 66332 0 -1 110976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_199_721
timestamp 1644511149
transform 1 0 67436 0 -1 110976
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_199_727
timestamp 1644511149
transform 1 0 67988 0 -1 110976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_199_729
timestamp 1644511149
transform 1 0 68172 0 -1 110976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_199_741
timestamp 1644511149
transform 1 0 69276 0 -1 110976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_199_753
timestamp 1644511149
transform 1 0 70380 0 -1 110976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_199_765
timestamp 1644511149
transform 1 0 71484 0 -1 110976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_199_777
timestamp 1644511149
transform 1 0 72588 0 -1 110976
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_199_783
timestamp 1644511149
transform 1 0 73140 0 -1 110976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_199_785
timestamp 1644511149
transform 1 0 73324 0 -1 110976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_199_797
timestamp 1644511149
transform 1 0 74428 0 -1 110976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_199_809
timestamp 1644511149
transform 1 0 75532 0 -1 110976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_199_821
timestamp 1644511149
transform 1 0 76636 0 -1 110976
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_199_829
timestamp 1644511149
transform 1 0 77372 0 -1 110976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_199_836
timestamp 1644511149
transform 1 0 78016 0 -1 110976
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_199_841
timestamp 1644511149
transform 1 0 78476 0 -1 110976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_200_3
timestamp 1644511149
transform 1 0 1380 0 1 110976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_200_15
timestamp 1644511149
transform 1 0 2484 0 1 110976
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_200_27
timestamp 1644511149
transform 1 0 3588 0 1 110976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_200_29
timestamp 1644511149
transform 1 0 3772 0 1 110976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_200_41
timestamp 1644511149
transform 1 0 4876 0 1 110976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_200_53
timestamp 1644511149
transform 1 0 5980 0 1 110976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_200_65
timestamp 1644511149
transform 1 0 7084 0 1 110976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_200_77
timestamp 1644511149
transform 1 0 8188 0 1 110976
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_200_83
timestamp 1644511149
transform 1 0 8740 0 1 110976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_200_85
timestamp 1644511149
transform 1 0 8924 0 1 110976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_200_97
timestamp 1644511149
transform 1 0 10028 0 1 110976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_200_109
timestamp 1644511149
transform 1 0 11132 0 1 110976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_200_121
timestamp 1644511149
transform 1 0 12236 0 1 110976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_200_133
timestamp 1644511149
transform 1 0 13340 0 1 110976
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_200_139
timestamp 1644511149
transform 1 0 13892 0 1 110976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_200_141
timestamp 1644511149
transform 1 0 14076 0 1 110976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_200_153
timestamp 1644511149
transform 1 0 15180 0 1 110976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_200_165
timestamp 1644511149
transform 1 0 16284 0 1 110976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_200_177
timestamp 1644511149
transform 1 0 17388 0 1 110976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_200_189
timestamp 1644511149
transform 1 0 18492 0 1 110976
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_200_195
timestamp 1644511149
transform 1 0 19044 0 1 110976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_200_197
timestamp 1644511149
transform 1 0 19228 0 1 110976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_200_209
timestamp 1644511149
transform 1 0 20332 0 1 110976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_200_221
timestamp 1644511149
transform 1 0 21436 0 1 110976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_200_233
timestamp 1644511149
transform 1 0 22540 0 1 110976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_200_245
timestamp 1644511149
transform 1 0 23644 0 1 110976
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_200_251
timestamp 1644511149
transform 1 0 24196 0 1 110976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_200_253
timestamp 1644511149
transform 1 0 24380 0 1 110976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_200_265
timestamp 1644511149
transform 1 0 25484 0 1 110976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_200_277
timestamp 1644511149
transform 1 0 26588 0 1 110976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_200_289
timestamp 1644511149
transform 1 0 27692 0 1 110976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_200_301
timestamp 1644511149
transform 1 0 28796 0 1 110976
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_200_307
timestamp 1644511149
transform 1 0 29348 0 1 110976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_200_309
timestamp 1644511149
transform 1 0 29532 0 1 110976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_200_321
timestamp 1644511149
transform 1 0 30636 0 1 110976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_200_333
timestamp 1644511149
transform 1 0 31740 0 1 110976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_200_345
timestamp 1644511149
transform 1 0 32844 0 1 110976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_200_357
timestamp 1644511149
transform 1 0 33948 0 1 110976
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_200_363
timestamp 1644511149
transform 1 0 34500 0 1 110976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_200_365
timestamp 1644511149
transform 1 0 34684 0 1 110976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_200_377
timestamp 1644511149
transform 1 0 35788 0 1 110976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_200_389
timestamp 1644511149
transform 1 0 36892 0 1 110976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_200_401
timestamp 1644511149
transform 1 0 37996 0 1 110976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_200_413
timestamp 1644511149
transform 1 0 39100 0 1 110976
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_200_419
timestamp 1644511149
transform 1 0 39652 0 1 110976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_200_421
timestamp 1644511149
transform 1 0 39836 0 1 110976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_200_433
timestamp 1644511149
transform 1 0 40940 0 1 110976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_200_445
timestamp 1644511149
transform 1 0 42044 0 1 110976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_200_457
timestamp 1644511149
transform 1 0 43148 0 1 110976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_200_469
timestamp 1644511149
transform 1 0 44252 0 1 110976
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_200_475
timestamp 1644511149
transform 1 0 44804 0 1 110976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_200_477
timestamp 1644511149
transform 1 0 44988 0 1 110976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_200_489
timestamp 1644511149
transform 1 0 46092 0 1 110976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_200_501
timestamp 1644511149
transform 1 0 47196 0 1 110976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_200_513
timestamp 1644511149
transform 1 0 48300 0 1 110976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_200_525
timestamp 1644511149
transform 1 0 49404 0 1 110976
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_200_531
timestamp 1644511149
transform 1 0 49956 0 1 110976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_200_533
timestamp 1644511149
transform 1 0 50140 0 1 110976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_200_545
timestamp 1644511149
transform 1 0 51244 0 1 110976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_200_557
timestamp 1644511149
transform 1 0 52348 0 1 110976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_200_569
timestamp 1644511149
transform 1 0 53452 0 1 110976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_200_581
timestamp 1644511149
transform 1 0 54556 0 1 110976
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_200_587
timestamp 1644511149
transform 1 0 55108 0 1 110976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_200_589
timestamp 1644511149
transform 1 0 55292 0 1 110976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_200_601
timestamp 1644511149
transform 1 0 56396 0 1 110976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_200_613
timestamp 1644511149
transform 1 0 57500 0 1 110976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_200_625
timestamp 1644511149
transform 1 0 58604 0 1 110976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_200_637
timestamp 1644511149
transform 1 0 59708 0 1 110976
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_200_643
timestamp 1644511149
transform 1 0 60260 0 1 110976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_200_645
timestamp 1644511149
transform 1 0 60444 0 1 110976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_200_657
timestamp 1644511149
transform 1 0 61548 0 1 110976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_200_669
timestamp 1644511149
transform 1 0 62652 0 1 110976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_200_681
timestamp 1644511149
transform 1 0 63756 0 1 110976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_200_693
timestamp 1644511149
transform 1 0 64860 0 1 110976
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_200_699
timestamp 1644511149
transform 1 0 65412 0 1 110976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_200_701
timestamp 1644511149
transform 1 0 65596 0 1 110976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_200_713
timestamp 1644511149
transform 1 0 66700 0 1 110976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_200_725
timestamp 1644511149
transform 1 0 67804 0 1 110976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_200_737
timestamp 1644511149
transform 1 0 68908 0 1 110976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_200_749
timestamp 1644511149
transform 1 0 70012 0 1 110976
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_200_755
timestamp 1644511149
transform 1 0 70564 0 1 110976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_200_757
timestamp 1644511149
transform 1 0 70748 0 1 110976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_200_769
timestamp 1644511149
transform 1 0 71852 0 1 110976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_200_781
timestamp 1644511149
transform 1 0 72956 0 1 110976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_200_793
timestamp 1644511149
transform 1 0 74060 0 1 110976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_200_805
timestamp 1644511149
transform 1 0 75164 0 1 110976
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_200_811
timestamp 1644511149
transform 1 0 75716 0 1 110976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_200_813
timestamp 1644511149
transform 1 0 75900 0 1 110976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_200_825
timestamp 1644511149
transform 1 0 77004 0 1 110976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_200_837
timestamp 1644511149
transform 1 0 78108 0 1 110976
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_200_841
timestamp 1644511149
transform 1 0 78476 0 1 110976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_201_3
timestamp 1644511149
transform 1 0 1380 0 -1 112064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_201_15
timestamp 1644511149
transform 1 0 2484 0 -1 112064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_201_27
timestamp 1644511149
transform 1 0 3588 0 -1 112064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_201_39
timestamp 1644511149
transform 1 0 4692 0 -1 112064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_201_51
timestamp 1644511149
transform 1 0 5796 0 -1 112064
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_201_55
timestamp 1644511149
transform 1 0 6164 0 -1 112064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_201_57
timestamp 1644511149
transform 1 0 6348 0 -1 112064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_201_69
timestamp 1644511149
transform 1 0 7452 0 -1 112064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_201_81
timestamp 1644511149
transform 1 0 8556 0 -1 112064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_201_93
timestamp 1644511149
transform 1 0 9660 0 -1 112064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_201_105
timestamp 1644511149
transform 1 0 10764 0 -1 112064
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_201_111
timestamp 1644511149
transform 1 0 11316 0 -1 112064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_201_113
timestamp 1644511149
transform 1 0 11500 0 -1 112064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_201_125
timestamp 1644511149
transform 1 0 12604 0 -1 112064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_201_137
timestamp 1644511149
transform 1 0 13708 0 -1 112064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_201_149
timestamp 1644511149
transform 1 0 14812 0 -1 112064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_201_161
timestamp 1644511149
transform 1 0 15916 0 -1 112064
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_201_167
timestamp 1644511149
transform 1 0 16468 0 -1 112064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_201_169
timestamp 1644511149
transform 1 0 16652 0 -1 112064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_201_181
timestamp 1644511149
transform 1 0 17756 0 -1 112064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_201_193
timestamp 1644511149
transform 1 0 18860 0 -1 112064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_201_205
timestamp 1644511149
transform 1 0 19964 0 -1 112064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_201_217
timestamp 1644511149
transform 1 0 21068 0 -1 112064
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_201_223
timestamp 1644511149
transform 1 0 21620 0 -1 112064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_201_225
timestamp 1644511149
transform 1 0 21804 0 -1 112064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_201_237
timestamp 1644511149
transform 1 0 22908 0 -1 112064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_201_249
timestamp 1644511149
transform 1 0 24012 0 -1 112064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_201_261
timestamp 1644511149
transform 1 0 25116 0 -1 112064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_201_273
timestamp 1644511149
transform 1 0 26220 0 -1 112064
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_201_279
timestamp 1644511149
transform 1 0 26772 0 -1 112064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_201_281
timestamp 1644511149
transform 1 0 26956 0 -1 112064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_201_293
timestamp 1644511149
transform 1 0 28060 0 -1 112064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_201_305
timestamp 1644511149
transform 1 0 29164 0 -1 112064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_201_317
timestamp 1644511149
transform 1 0 30268 0 -1 112064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_201_329
timestamp 1644511149
transform 1 0 31372 0 -1 112064
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_201_335
timestamp 1644511149
transform 1 0 31924 0 -1 112064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_201_337
timestamp 1644511149
transform 1 0 32108 0 -1 112064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_201_349
timestamp 1644511149
transform 1 0 33212 0 -1 112064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_201_361
timestamp 1644511149
transform 1 0 34316 0 -1 112064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_201_373
timestamp 1644511149
transform 1 0 35420 0 -1 112064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_201_385
timestamp 1644511149
transform 1 0 36524 0 -1 112064
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_201_391
timestamp 1644511149
transform 1 0 37076 0 -1 112064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_201_393
timestamp 1644511149
transform 1 0 37260 0 -1 112064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_201_405
timestamp 1644511149
transform 1 0 38364 0 -1 112064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_201_417
timestamp 1644511149
transform 1 0 39468 0 -1 112064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_201_429
timestamp 1644511149
transform 1 0 40572 0 -1 112064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_201_441
timestamp 1644511149
transform 1 0 41676 0 -1 112064
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_201_447
timestamp 1644511149
transform 1 0 42228 0 -1 112064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_201_449
timestamp 1644511149
transform 1 0 42412 0 -1 112064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_201_461
timestamp 1644511149
transform 1 0 43516 0 -1 112064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_201_473
timestamp 1644511149
transform 1 0 44620 0 -1 112064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_201_485
timestamp 1644511149
transform 1 0 45724 0 -1 112064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_201_497
timestamp 1644511149
transform 1 0 46828 0 -1 112064
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_201_503
timestamp 1644511149
transform 1 0 47380 0 -1 112064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_201_505
timestamp 1644511149
transform 1 0 47564 0 -1 112064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_201_517
timestamp 1644511149
transform 1 0 48668 0 -1 112064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_201_529
timestamp 1644511149
transform 1 0 49772 0 -1 112064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_201_541
timestamp 1644511149
transform 1 0 50876 0 -1 112064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_201_553
timestamp 1644511149
transform 1 0 51980 0 -1 112064
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_201_559
timestamp 1644511149
transform 1 0 52532 0 -1 112064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_201_561
timestamp 1644511149
transform 1 0 52716 0 -1 112064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_201_573
timestamp 1644511149
transform 1 0 53820 0 -1 112064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_201_585
timestamp 1644511149
transform 1 0 54924 0 -1 112064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_201_597
timestamp 1644511149
transform 1 0 56028 0 -1 112064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_201_609
timestamp 1644511149
transform 1 0 57132 0 -1 112064
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_201_615
timestamp 1644511149
transform 1 0 57684 0 -1 112064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_201_617
timestamp 1644511149
transform 1 0 57868 0 -1 112064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_201_629
timestamp 1644511149
transform 1 0 58972 0 -1 112064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_201_641
timestamp 1644511149
transform 1 0 60076 0 -1 112064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_201_653
timestamp 1644511149
transform 1 0 61180 0 -1 112064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_201_665
timestamp 1644511149
transform 1 0 62284 0 -1 112064
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_201_671
timestamp 1644511149
transform 1 0 62836 0 -1 112064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_201_673
timestamp 1644511149
transform 1 0 63020 0 -1 112064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_201_685
timestamp 1644511149
transform 1 0 64124 0 -1 112064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_201_697
timestamp 1644511149
transform 1 0 65228 0 -1 112064
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_201_709
timestamp 1644511149
transform 1 0 66332 0 -1 112064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_201_714
timestamp 1644511149
transform 1 0 66792 0 -1 112064
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_201_726
timestamp 1644511149
transform 1 0 67896 0 -1 112064
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_201_729
timestamp 1644511149
transform 1 0 68172 0 -1 112064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_201_741
timestamp 1644511149
transform 1 0 69276 0 -1 112064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_201_753
timestamp 1644511149
transform 1 0 70380 0 -1 112064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_201_765
timestamp 1644511149
transform 1 0 71484 0 -1 112064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_201_777
timestamp 1644511149
transform 1 0 72588 0 -1 112064
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_201_783
timestamp 1644511149
transform 1 0 73140 0 -1 112064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_201_785
timestamp 1644511149
transform 1 0 73324 0 -1 112064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_201_797
timestamp 1644511149
transform 1 0 74428 0 -1 112064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_201_809
timestamp 1644511149
transform 1 0 75532 0 -1 112064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_201_821
timestamp 1644511149
transform 1 0 76636 0 -1 112064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_201_833
timestamp 1644511149
transform 1 0 77740 0 -1 112064
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_201_839
timestamp 1644511149
transform 1 0 78292 0 -1 112064
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_201_841
timestamp 1644511149
transform 1 0 78476 0 -1 112064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_202_3
timestamp 1644511149
transform 1 0 1380 0 1 112064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_202_15
timestamp 1644511149
transform 1 0 2484 0 1 112064
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_202_27
timestamp 1644511149
transform 1 0 3588 0 1 112064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_202_29
timestamp 1644511149
transform 1 0 3772 0 1 112064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_202_41
timestamp 1644511149
transform 1 0 4876 0 1 112064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_202_53
timestamp 1644511149
transform 1 0 5980 0 1 112064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_202_65
timestamp 1644511149
transform 1 0 7084 0 1 112064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_202_77
timestamp 1644511149
transform 1 0 8188 0 1 112064
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_202_83
timestamp 1644511149
transform 1 0 8740 0 1 112064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_202_85
timestamp 1644511149
transform 1 0 8924 0 1 112064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_202_97
timestamp 1644511149
transform 1 0 10028 0 1 112064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_202_109
timestamp 1644511149
transform 1 0 11132 0 1 112064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_202_121
timestamp 1644511149
transform 1 0 12236 0 1 112064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_202_133
timestamp 1644511149
transform 1 0 13340 0 1 112064
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_202_139
timestamp 1644511149
transform 1 0 13892 0 1 112064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_202_141
timestamp 1644511149
transform 1 0 14076 0 1 112064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_202_153
timestamp 1644511149
transform 1 0 15180 0 1 112064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_202_165
timestamp 1644511149
transform 1 0 16284 0 1 112064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_202_177
timestamp 1644511149
transform 1 0 17388 0 1 112064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_202_189
timestamp 1644511149
transform 1 0 18492 0 1 112064
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_202_195
timestamp 1644511149
transform 1 0 19044 0 1 112064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_202_197
timestamp 1644511149
transform 1 0 19228 0 1 112064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_202_209
timestamp 1644511149
transform 1 0 20332 0 1 112064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_202_221
timestamp 1644511149
transform 1 0 21436 0 1 112064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_202_233
timestamp 1644511149
transform 1 0 22540 0 1 112064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_202_245
timestamp 1644511149
transform 1 0 23644 0 1 112064
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_202_251
timestamp 1644511149
transform 1 0 24196 0 1 112064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_202_253
timestamp 1644511149
transform 1 0 24380 0 1 112064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_202_265
timestamp 1644511149
transform 1 0 25484 0 1 112064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_202_277
timestamp 1644511149
transform 1 0 26588 0 1 112064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_202_289
timestamp 1644511149
transform 1 0 27692 0 1 112064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_202_301
timestamp 1644511149
transform 1 0 28796 0 1 112064
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_202_307
timestamp 1644511149
transform 1 0 29348 0 1 112064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_202_309
timestamp 1644511149
transform 1 0 29532 0 1 112064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_202_321
timestamp 1644511149
transform 1 0 30636 0 1 112064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_202_333
timestamp 1644511149
transform 1 0 31740 0 1 112064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_202_345
timestamp 1644511149
transform 1 0 32844 0 1 112064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_202_357
timestamp 1644511149
transform 1 0 33948 0 1 112064
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_202_363
timestamp 1644511149
transform 1 0 34500 0 1 112064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_202_365
timestamp 1644511149
transform 1 0 34684 0 1 112064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_202_377
timestamp 1644511149
transform 1 0 35788 0 1 112064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_202_389
timestamp 1644511149
transform 1 0 36892 0 1 112064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_202_401
timestamp 1644511149
transform 1 0 37996 0 1 112064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_202_413
timestamp 1644511149
transform 1 0 39100 0 1 112064
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_202_419
timestamp 1644511149
transform 1 0 39652 0 1 112064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_202_421
timestamp 1644511149
transform 1 0 39836 0 1 112064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_202_433
timestamp 1644511149
transform 1 0 40940 0 1 112064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_202_445
timestamp 1644511149
transform 1 0 42044 0 1 112064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_202_457
timestamp 1644511149
transform 1 0 43148 0 1 112064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_202_469
timestamp 1644511149
transform 1 0 44252 0 1 112064
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_202_475
timestamp 1644511149
transform 1 0 44804 0 1 112064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_202_477
timestamp 1644511149
transform 1 0 44988 0 1 112064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_202_489
timestamp 1644511149
transform 1 0 46092 0 1 112064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_202_501
timestamp 1644511149
transform 1 0 47196 0 1 112064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_202_513
timestamp 1644511149
transform 1 0 48300 0 1 112064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_202_525
timestamp 1644511149
transform 1 0 49404 0 1 112064
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_202_531
timestamp 1644511149
transform 1 0 49956 0 1 112064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_202_533
timestamp 1644511149
transform 1 0 50140 0 1 112064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_202_545
timestamp 1644511149
transform 1 0 51244 0 1 112064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_202_557
timestamp 1644511149
transform 1 0 52348 0 1 112064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_202_569
timestamp 1644511149
transform 1 0 53452 0 1 112064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_202_581
timestamp 1644511149
transform 1 0 54556 0 1 112064
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_202_587
timestamp 1644511149
transform 1 0 55108 0 1 112064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_202_589
timestamp 1644511149
transform 1 0 55292 0 1 112064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_202_601
timestamp 1644511149
transform 1 0 56396 0 1 112064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_202_613
timestamp 1644511149
transform 1 0 57500 0 1 112064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_202_625
timestamp 1644511149
transform 1 0 58604 0 1 112064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_202_637
timestamp 1644511149
transform 1 0 59708 0 1 112064
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_202_643
timestamp 1644511149
transform 1 0 60260 0 1 112064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_202_645
timestamp 1644511149
transform 1 0 60444 0 1 112064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_202_657
timestamp 1644511149
transform 1 0 61548 0 1 112064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_202_669
timestamp 1644511149
transform 1 0 62652 0 1 112064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_202_681
timestamp 1644511149
transform 1 0 63756 0 1 112064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_202_693
timestamp 1644511149
transform 1 0 64860 0 1 112064
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_202_699
timestamp 1644511149
transform 1 0 65412 0 1 112064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_202_701
timestamp 1644511149
transform 1 0 65596 0 1 112064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_202_713
timestamp 1644511149
transform 1 0 66700 0 1 112064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_202_725
timestamp 1644511149
transform 1 0 67804 0 1 112064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_202_737
timestamp 1644511149
transform 1 0 68908 0 1 112064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_202_749
timestamp 1644511149
transform 1 0 70012 0 1 112064
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_202_755
timestamp 1644511149
transform 1 0 70564 0 1 112064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_202_757
timestamp 1644511149
transform 1 0 70748 0 1 112064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_202_769
timestamp 1644511149
transform 1 0 71852 0 1 112064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_202_781
timestamp 1644511149
transform 1 0 72956 0 1 112064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_202_793
timestamp 1644511149
transform 1 0 74060 0 1 112064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_202_805
timestamp 1644511149
transform 1 0 75164 0 1 112064
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_202_811
timestamp 1644511149
transform 1 0 75716 0 1 112064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_202_813
timestamp 1644511149
transform 1 0 75900 0 1 112064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_202_825
timestamp 1644511149
transform 1 0 77004 0 1 112064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_202_837
timestamp 1644511149
transform 1 0 78108 0 1 112064
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_202_841
timestamp 1644511149
transform 1 0 78476 0 1 112064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_203_3
timestamp 1644511149
transform 1 0 1380 0 -1 113152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_203_15
timestamp 1644511149
transform 1 0 2484 0 -1 113152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_203_27
timestamp 1644511149
transform 1 0 3588 0 -1 113152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_203_39
timestamp 1644511149
transform 1 0 4692 0 -1 113152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_203_51
timestamp 1644511149
transform 1 0 5796 0 -1 113152
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_203_55
timestamp 1644511149
transform 1 0 6164 0 -1 113152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_203_57
timestamp 1644511149
transform 1 0 6348 0 -1 113152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_203_69
timestamp 1644511149
transform 1 0 7452 0 -1 113152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_203_81
timestamp 1644511149
transform 1 0 8556 0 -1 113152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_203_93
timestamp 1644511149
transform 1 0 9660 0 -1 113152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_203_105
timestamp 1644511149
transform 1 0 10764 0 -1 113152
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_203_111
timestamp 1644511149
transform 1 0 11316 0 -1 113152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_203_113
timestamp 1644511149
transform 1 0 11500 0 -1 113152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_203_125
timestamp 1644511149
transform 1 0 12604 0 -1 113152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_203_137
timestamp 1644511149
transform 1 0 13708 0 -1 113152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_203_149
timestamp 1644511149
transform 1 0 14812 0 -1 113152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_203_161
timestamp 1644511149
transform 1 0 15916 0 -1 113152
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_203_167
timestamp 1644511149
transform 1 0 16468 0 -1 113152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_203_169
timestamp 1644511149
transform 1 0 16652 0 -1 113152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_203_181
timestamp 1644511149
transform 1 0 17756 0 -1 113152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_203_193
timestamp 1644511149
transform 1 0 18860 0 -1 113152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_203_205
timestamp 1644511149
transform 1 0 19964 0 -1 113152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_203_217
timestamp 1644511149
transform 1 0 21068 0 -1 113152
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_203_223
timestamp 1644511149
transform 1 0 21620 0 -1 113152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_203_225
timestamp 1644511149
transform 1 0 21804 0 -1 113152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_203_237
timestamp 1644511149
transform 1 0 22908 0 -1 113152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_203_249
timestamp 1644511149
transform 1 0 24012 0 -1 113152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_203_261
timestamp 1644511149
transform 1 0 25116 0 -1 113152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_203_273
timestamp 1644511149
transform 1 0 26220 0 -1 113152
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_203_279
timestamp 1644511149
transform 1 0 26772 0 -1 113152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_203_281
timestamp 1644511149
transform 1 0 26956 0 -1 113152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_203_293
timestamp 1644511149
transform 1 0 28060 0 -1 113152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_203_305
timestamp 1644511149
transform 1 0 29164 0 -1 113152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_203_317
timestamp 1644511149
transform 1 0 30268 0 -1 113152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_203_329
timestamp 1644511149
transform 1 0 31372 0 -1 113152
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_203_335
timestamp 1644511149
transform 1 0 31924 0 -1 113152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_203_337
timestamp 1644511149
transform 1 0 32108 0 -1 113152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_203_349
timestamp 1644511149
transform 1 0 33212 0 -1 113152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_203_361
timestamp 1644511149
transform 1 0 34316 0 -1 113152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_203_373
timestamp 1644511149
transform 1 0 35420 0 -1 113152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_203_385
timestamp 1644511149
transform 1 0 36524 0 -1 113152
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_203_391
timestamp 1644511149
transform 1 0 37076 0 -1 113152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_203_393
timestamp 1644511149
transform 1 0 37260 0 -1 113152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_203_405
timestamp 1644511149
transform 1 0 38364 0 -1 113152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_203_417
timestamp 1644511149
transform 1 0 39468 0 -1 113152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_203_429
timestamp 1644511149
transform 1 0 40572 0 -1 113152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_203_441
timestamp 1644511149
transform 1 0 41676 0 -1 113152
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_203_447
timestamp 1644511149
transform 1 0 42228 0 -1 113152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_203_449
timestamp 1644511149
transform 1 0 42412 0 -1 113152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_203_461
timestamp 1644511149
transform 1 0 43516 0 -1 113152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_203_473
timestamp 1644511149
transform 1 0 44620 0 -1 113152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_203_485
timestamp 1644511149
transform 1 0 45724 0 -1 113152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_203_497
timestamp 1644511149
transform 1 0 46828 0 -1 113152
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_203_503
timestamp 1644511149
transform 1 0 47380 0 -1 113152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_203_505
timestamp 1644511149
transform 1 0 47564 0 -1 113152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_203_517
timestamp 1644511149
transform 1 0 48668 0 -1 113152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_203_529
timestamp 1644511149
transform 1 0 49772 0 -1 113152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_203_541
timestamp 1644511149
transform 1 0 50876 0 -1 113152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_203_553
timestamp 1644511149
transform 1 0 51980 0 -1 113152
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_203_559
timestamp 1644511149
transform 1 0 52532 0 -1 113152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_203_561
timestamp 1644511149
transform 1 0 52716 0 -1 113152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_203_573
timestamp 1644511149
transform 1 0 53820 0 -1 113152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_203_585
timestamp 1644511149
transform 1 0 54924 0 -1 113152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_203_597
timestamp 1644511149
transform 1 0 56028 0 -1 113152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_203_609
timestamp 1644511149
transform 1 0 57132 0 -1 113152
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_203_615
timestamp 1644511149
transform 1 0 57684 0 -1 113152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_203_617
timestamp 1644511149
transform 1 0 57868 0 -1 113152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_203_629
timestamp 1644511149
transform 1 0 58972 0 -1 113152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_203_641
timestamp 1644511149
transform 1 0 60076 0 -1 113152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_203_653
timestamp 1644511149
transform 1 0 61180 0 -1 113152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_203_665
timestamp 1644511149
transform 1 0 62284 0 -1 113152
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_203_671
timestamp 1644511149
transform 1 0 62836 0 -1 113152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_203_673
timestamp 1644511149
transform 1 0 63020 0 -1 113152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_203_685
timestamp 1644511149
transform 1 0 64124 0 -1 113152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_203_697
timestamp 1644511149
transform 1 0 65228 0 -1 113152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_203_709
timestamp 1644511149
transform 1 0 66332 0 -1 113152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_203_721
timestamp 1644511149
transform 1 0 67436 0 -1 113152
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_203_727
timestamp 1644511149
transform 1 0 67988 0 -1 113152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_203_729
timestamp 1644511149
transform 1 0 68172 0 -1 113152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_203_741
timestamp 1644511149
transform 1 0 69276 0 -1 113152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_203_753
timestamp 1644511149
transform 1 0 70380 0 -1 113152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_203_765
timestamp 1644511149
transform 1 0 71484 0 -1 113152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_203_777
timestamp 1644511149
transform 1 0 72588 0 -1 113152
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_203_783
timestamp 1644511149
transform 1 0 73140 0 -1 113152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_203_785
timestamp 1644511149
transform 1 0 73324 0 -1 113152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_203_797
timestamp 1644511149
transform 1 0 74428 0 -1 113152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_203_809
timestamp 1644511149
transform 1 0 75532 0 -1 113152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_203_821
timestamp 1644511149
transform 1 0 76636 0 -1 113152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_203_833
timestamp 1644511149
transform 1 0 77740 0 -1 113152
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_203_839
timestamp 1644511149
transform 1 0 78292 0 -1 113152
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_203_841
timestamp 1644511149
transform 1 0 78476 0 -1 113152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_204_7
timestamp 1644511149
transform 1 0 1748 0 1 113152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_204_19
timestamp 1644511149
transform 1 0 2852 0 1 113152
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_204_27
timestamp 1644511149
transform 1 0 3588 0 1 113152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_204_29
timestamp 1644511149
transform 1 0 3772 0 1 113152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_204_41
timestamp 1644511149
transform 1 0 4876 0 1 113152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_204_53
timestamp 1644511149
transform 1 0 5980 0 1 113152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_204_65
timestamp 1644511149
transform 1 0 7084 0 1 113152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_204_77
timestamp 1644511149
transform 1 0 8188 0 1 113152
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_204_83
timestamp 1644511149
transform 1 0 8740 0 1 113152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_204_85
timestamp 1644511149
transform 1 0 8924 0 1 113152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_204_97
timestamp 1644511149
transform 1 0 10028 0 1 113152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_204_109
timestamp 1644511149
transform 1 0 11132 0 1 113152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_204_121
timestamp 1644511149
transform 1 0 12236 0 1 113152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_204_133
timestamp 1644511149
transform 1 0 13340 0 1 113152
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_204_139
timestamp 1644511149
transform 1 0 13892 0 1 113152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_204_141
timestamp 1644511149
transform 1 0 14076 0 1 113152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_204_153
timestamp 1644511149
transform 1 0 15180 0 1 113152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_204_165
timestamp 1644511149
transform 1 0 16284 0 1 113152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_204_177
timestamp 1644511149
transform 1 0 17388 0 1 113152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_204_189
timestamp 1644511149
transform 1 0 18492 0 1 113152
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_204_195
timestamp 1644511149
transform 1 0 19044 0 1 113152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_204_197
timestamp 1644511149
transform 1 0 19228 0 1 113152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_204_209
timestamp 1644511149
transform 1 0 20332 0 1 113152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_204_221
timestamp 1644511149
transform 1 0 21436 0 1 113152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_204_233
timestamp 1644511149
transform 1 0 22540 0 1 113152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_204_245
timestamp 1644511149
transform 1 0 23644 0 1 113152
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_204_251
timestamp 1644511149
transform 1 0 24196 0 1 113152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_204_253
timestamp 1644511149
transform 1 0 24380 0 1 113152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_204_265
timestamp 1644511149
transform 1 0 25484 0 1 113152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_204_277
timestamp 1644511149
transform 1 0 26588 0 1 113152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_204_289
timestamp 1644511149
transform 1 0 27692 0 1 113152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_204_301
timestamp 1644511149
transform 1 0 28796 0 1 113152
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_204_307
timestamp 1644511149
transform 1 0 29348 0 1 113152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_204_309
timestamp 1644511149
transform 1 0 29532 0 1 113152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_204_321
timestamp 1644511149
transform 1 0 30636 0 1 113152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_204_333
timestamp 1644511149
transform 1 0 31740 0 1 113152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_204_345
timestamp 1644511149
transform 1 0 32844 0 1 113152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_204_357
timestamp 1644511149
transform 1 0 33948 0 1 113152
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_204_363
timestamp 1644511149
transform 1 0 34500 0 1 113152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_204_365
timestamp 1644511149
transform 1 0 34684 0 1 113152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_204_377
timestamp 1644511149
transform 1 0 35788 0 1 113152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_204_389
timestamp 1644511149
transform 1 0 36892 0 1 113152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_204_401
timestamp 1644511149
transform 1 0 37996 0 1 113152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_204_413
timestamp 1644511149
transform 1 0 39100 0 1 113152
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_204_419
timestamp 1644511149
transform 1 0 39652 0 1 113152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_204_421
timestamp 1644511149
transform 1 0 39836 0 1 113152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_204_433
timestamp 1644511149
transform 1 0 40940 0 1 113152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_204_445
timestamp 1644511149
transform 1 0 42044 0 1 113152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_204_457
timestamp 1644511149
transform 1 0 43148 0 1 113152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_204_469
timestamp 1644511149
transform 1 0 44252 0 1 113152
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_204_475
timestamp 1644511149
transform 1 0 44804 0 1 113152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_204_477
timestamp 1644511149
transform 1 0 44988 0 1 113152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_204_489
timestamp 1644511149
transform 1 0 46092 0 1 113152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_204_501
timestamp 1644511149
transform 1 0 47196 0 1 113152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_204_513
timestamp 1644511149
transform 1 0 48300 0 1 113152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_204_525
timestamp 1644511149
transform 1 0 49404 0 1 113152
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_204_531
timestamp 1644511149
transform 1 0 49956 0 1 113152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_204_533
timestamp 1644511149
transform 1 0 50140 0 1 113152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_204_545
timestamp 1644511149
transform 1 0 51244 0 1 113152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_204_557
timestamp 1644511149
transform 1 0 52348 0 1 113152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_204_569
timestamp 1644511149
transform 1 0 53452 0 1 113152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_204_581
timestamp 1644511149
transform 1 0 54556 0 1 113152
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_204_587
timestamp 1644511149
transform 1 0 55108 0 1 113152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_204_589
timestamp 1644511149
transform 1 0 55292 0 1 113152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_204_601
timestamp 1644511149
transform 1 0 56396 0 1 113152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_204_613
timestamp 1644511149
transform 1 0 57500 0 1 113152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_204_625
timestamp 1644511149
transform 1 0 58604 0 1 113152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_204_637
timestamp 1644511149
transform 1 0 59708 0 1 113152
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_204_643
timestamp 1644511149
transform 1 0 60260 0 1 113152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_204_645
timestamp 1644511149
transform 1 0 60444 0 1 113152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_204_657
timestamp 1644511149
transform 1 0 61548 0 1 113152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_204_669
timestamp 1644511149
transform 1 0 62652 0 1 113152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_204_681
timestamp 1644511149
transform 1 0 63756 0 1 113152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_204_693
timestamp 1644511149
transform 1 0 64860 0 1 113152
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_204_699
timestamp 1644511149
transform 1 0 65412 0 1 113152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_204_701
timestamp 1644511149
transform 1 0 65596 0 1 113152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_204_713
timestamp 1644511149
transform 1 0 66700 0 1 113152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_204_725
timestamp 1644511149
transform 1 0 67804 0 1 113152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_204_737
timestamp 1644511149
transform 1 0 68908 0 1 113152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_204_749
timestamp 1644511149
transform 1 0 70012 0 1 113152
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_204_755
timestamp 1644511149
transform 1 0 70564 0 1 113152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_204_757
timestamp 1644511149
transform 1 0 70748 0 1 113152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_204_769
timestamp 1644511149
transform 1 0 71852 0 1 113152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_204_781
timestamp 1644511149
transform 1 0 72956 0 1 113152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_204_793
timestamp 1644511149
transform 1 0 74060 0 1 113152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_204_805
timestamp 1644511149
transform 1 0 75164 0 1 113152
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_204_811
timestamp 1644511149
transform 1 0 75716 0 1 113152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_204_813
timestamp 1644511149
transform 1 0 75900 0 1 113152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_204_825
timestamp 1644511149
transform 1 0 77004 0 1 113152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_204_837
timestamp 1644511149
transform 1 0 78108 0 1 113152
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_204_841
timestamp 1644511149
transform 1 0 78476 0 1 113152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_205_3
timestamp 1644511149
transform 1 0 1380 0 -1 114240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_205_15
timestamp 1644511149
transform 1 0 2484 0 -1 114240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_205_27
timestamp 1644511149
transform 1 0 3588 0 -1 114240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_205_39
timestamp 1644511149
transform 1 0 4692 0 -1 114240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_205_51
timestamp 1644511149
transform 1 0 5796 0 -1 114240
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_205_55
timestamp 1644511149
transform 1 0 6164 0 -1 114240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_205_57
timestamp 1644511149
transform 1 0 6348 0 -1 114240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_205_69
timestamp 1644511149
transform 1 0 7452 0 -1 114240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_205_81
timestamp 1644511149
transform 1 0 8556 0 -1 114240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_205_93
timestamp 1644511149
transform 1 0 9660 0 -1 114240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_205_105
timestamp 1644511149
transform 1 0 10764 0 -1 114240
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_205_111
timestamp 1644511149
transform 1 0 11316 0 -1 114240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_205_113
timestamp 1644511149
transform 1 0 11500 0 -1 114240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_205_125
timestamp 1644511149
transform 1 0 12604 0 -1 114240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_205_137
timestamp 1644511149
transform 1 0 13708 0 -1 114240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_205_149
timestamp 1644511149
transform 1 0 14812 0 -1 114240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_205_161
timestamp 1644511149
transform 1 0 15916 0 -1 114240
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_205_167
timestamp 1644511149
transform 1 0 16468 0 -1 114240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_205_169
timestamp 1644511149
transform 1 0 16652 0 -1 114240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_205_181
timestamp 1644511149
transform 1 0 17756 0 -1 114240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_205_193
timestamp 1644511149
transform 1 0 18860 0 -1 114240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_205_205
timestamp 1644511149
transform 1 0 19964 0 -1 114240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_205_217
timestamp 1644511149
transform 1 0 21068 0 -1 114240
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_205_223
timestamp 1644511149
transform 1 0 21620 0 -1 114240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_205_225
timestamp 1644511149
transform 1 0 21804 0 -1 114240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_205_237
timestamp 1644511149
transform 1 0 22908 0 -1 114240
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_205_249
timestamp 1644511149
transform 1 0 24012 0 -1 114240
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_205_254
timestamp 1644511149
transform 1 0 24472 0 -1 114240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_205_266
timestamp 1644511149
transform 1 0 25576 0 -1 114240
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_205_278
timestamp 1644511149
transform 1 0 26680 0 -1 114240
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_205_281
timestamp 1644511149
transform 1 0 26956 0 -1 114240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_205_293
timestamp 1644511149
transform 1 0 28060 0 -1 114240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_205_305
timestamp 1644511149
transform 1 0 29164 0 -1 114240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_205_317
timestamp 1644511149
transform 1 0 30268 0 -1 114240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_205_329
timestamp 1644511149
transform 1 0 31372 0 -1 114240
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_205_335
timestamp 1644511149
transform 1 0 31924 0 -1 114240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_205_337
timestamp 1644511149
transform 1 0 32108 0 -1 114240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_205_349
timestamp 1644511149
transform 1 0 33212 0 -1 114240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_205_361
timestamp 1644511149
transform 1 0 34316 0 -1 114240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_205_373
timestamp 1644511149
transform 1 0 35420 0 -1 114240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_205_385
timestamp 1644511149
transform 1 0 36524 0 -1 114240
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_205_391
timestamp 1644511149
transform 1 0 37076 0 -1 114240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_205_393
timestamp 1644511149
transform 1 0 37260 0 -1 114240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_205_405
timestamp 1644511149
transform 1 0 38364 0 -1 114240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_205_417
timestamp 1644511149
transform 1 0 39468 0 -1 114240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_205_429
timestamp 1644511149
transform 1 0 40572 0 -1 114240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_205_441
timestamp 1644511149
transform 1 0 41676 0 -1 114240
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_205_447
timestamp 1644511149
transform 1 0 42228 0 -1 114240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_205_449
timestamp 1644511149
transform 1 0 42412 0 -1 114240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_205_461
timestamp 1644511149
transform 1 0 43516 0 -1 114240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_205_473
timestamp 1644511149
transform 1 0 44620 0 -1 114240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_205_485
timestamp 1644511149
transform 1 0 45724 0 -1 114240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_205_497
timestamp 1644511149
transform 1 0 46828 0 -1 114240
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_205_503
timestamp 1644511149
transform 1 0 47380 0 -1 114240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_205_505
timestamp 1644511149
transform 1 0 47564 0 -1 114240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_205_517
timestamp 1644511149
transform 1 0 48668 0 -1 114240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_205_529
timestamp 1644511149
transform 1 0 49772 0 -1 114240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_205_541
timestamp 1644511149
transform 1 0 50876 0 -1 114240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_205_553
timestamp 1644511149
transform 1 0 51980 0 -1 114240
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_205_559
timestamp 1644511149
transform 1 0 52532 0 -1 114240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_205_561
timestamp 1644511149
transform 1 0 52716 0 -1 114240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_205_573
timestamp 1644511149
transform 1 0 53820 0 -1 114240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_205_585
timestamp 1644511149
transform 1 0 54924 0 -1 114240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_205_597
timestamp 1644511149
transform 1 0 56028 0 -1 114240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_205_609
timestamp 1644511149
transform 1 0 57132 0 -1 114240
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_205_615
timestamp 1644511149
transform 1 0 57684 0 -1 114240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_205_617
timestamp 1644511149
transform 1 0 57868 0 -1 114240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_205_629
timestamp 1644511149
transform 1 0 58972 0 -1 114240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_205_641
timestamp 1644511149
transform 1 0 60076 0 -1 114240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_205_653
timestamp 1644511149
transform 1 0 61180 0 -1 114240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_205_665
timestamp 1644511149
transform 1 0 62284 0 -1 114240
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_205_671
timestamp 1644511149
transform 1 0 62836 0 -1 114240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_205_673
timestamp 1644511149
transform 1 0 63020 0 -1 114240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_205_685
timestamp 1644511149
transform 1 0 64124 0 -1 114240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_205_697
timestamp 1644511149
transform 1 0 65228 0 -1 114240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_205_709
timestamp 1644511149
transform 1 0 66332 0 -1 114240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_205_721
timestamp 1644511149
transform 1 0 67436 0 -1 114240
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_205_727
timestamp 1644511149
transform 1 0 67988 0 -1 114240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_205_729
timestamp 1644511149
transform 1 0 68172 0 -1 114240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_205_741
timestamp 1644511149
transform 1 0 69276 0 -1 114240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_205_753
timestamp 1644511149
transform 1 0 70380 0 -1 114240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_205_765
timestamp 1644511149
transform 1 0 71484 0 -1 114240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_205_777
timestamp 1644511149
transform 1 0 72588 0 -1 114240
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_205_783
timestamp 1644511149
transform 1 0 73140 0 -1 114240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_205_785
timestamp 1644511149
transform 1 0 73324 0 -1 114240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_205_797
timestamp 1644511149
transform 1 0 74428 0 -1 114240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_205_809
timestamp 1644511149
transform 1 0 75532 0 -1 114240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_205_821
timestamp 1644511149
transform 1 0 76636 0 -1 114240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_205_833
timestamp 1644511149
transform 1 0 77740 0 -1 114240
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_205_839
timestamp 1644511149
transform 1 0 78292 0 -1 114240
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_205_841
timestamp 1644511149
transform 1 0 78476 0 -1 114240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_206_3
timestamp 1644511149
transform 1 0 1380 0 1 114240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_206_15
timestamp 1644511149
transform 1 0 2484 0 1 114240
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_206_27
timestamp 1644511149
transform 1 0 3588 0 1 114240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_206_29
timestamp 1644511149
transform 1 0 3772 0 1 114240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_206_41
timestamp 1644511149
transform 1 0 4876 0 1 114240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_206_53
timestamp 1644511149
transform 1 0 5980 0 1 114240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_206_65
timestamp 1644511149
transform 1 0 7084 0 1 114240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_206_77
timestamp 1644511149
transform 1 0 8188 0 1 114240
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_206_83
timestamp 1644511149
transform 1 0 8740 0 1 114240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_206_85
timestamp 1644511149
transform 1 0 8924 0 1 114240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_206_97
timestamp 1644511149
transform 1 0 10028 0 1 114240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_206_109
timestamp 1644511149
transform 1 0 11132 0 1 114240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_206_121
timestamp 1644511149
transform 1 0 12236 0 1 114240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_206_133
timestamp 1644511149
transform 1 0 13340 0 1 114240
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_206_139
timestamp 1644511149
transform 1 0 13892 0 1 114240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_206_141
timestamp 1644511149
transform 1 0 14076 0 1 114240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_206_153
timestamp 1644511149
transform 1 0 15180 0 1 114240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_206_165
timestamp 1644511149
transform 1 0 16284 0 1 114240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_206_177
timestamp 1644511149
transform 1 0 17388 0 1 114240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_206_189
timestamp 1644511149
transform 1 0 18492 0 1 114240
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_206_195
timestamp 1644511149
transform 1 0 19044 0 1 114240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_206_197
timestamp 1644511149
transform 1 0 19228 0 1 114240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_206_209
timestamp 1644511149
transform 1 0 20332 0 1 114240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_206_221
timestamp 1644511149
transform 1 0 21436 0 1 114240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_206_233
timestamp 1644511149
transform 1 0 22540 0 1 114240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_206_245
timestamp 1644511149
transform 1 0 23644 0 1 114240
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_206_251
timestamp 1644511149
transform 1 0 24196 0 1 114240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_206_253
timestamp 1644511149
transform 1 0 24380 0 1 114240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_206_265
timestamp 1644511149
transform 1 0 25484 0 1 114240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_206_277
timestamp 1644511149
transform 1 0 26588 0 1 114240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_206_289
timestamp 1644511149
transform 1 0 27692 0 1 114240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_206_301
timestamp 1644511149
transform 1 0 28796 0 1 114240
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_206_307
timestamp 1644511149
transform 1 0 29348 0 1 114240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_206_309
timestamp 1644511149
transform 1 0 29532 0 1 114240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_206_321
timestamp 1644511149
transform 1 0 30636 0 1 114240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_206_333
timestamp 1644511149
transform 1 0 31740 0 1 114240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_206_345
timestamp 1644511149
transform 1 0 32844 0 1 114240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_206_357
timestamp 1644511149
transform 1 0 33948 0 1 114240
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_206_363
timestamp 1644511149
transform 1 0 34500 0 1 114240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_206_365
timestamp 1644511149
transform 1 0 34684 0 1 114240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_206_377
timestamp 1644511149
transform 1 0 35788 0 1 114240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_206_389
timestamp 1644511149
transform 1 0 36892 0 1 114240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_206_401
timestamp 1644511149
transform 1 0 37996 0 1 114240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_206_413
timestamp 1644511149
transform 1 0 39100 0 1 114240
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_206_419
timestamp 1644511149
transform 1 0 39652 0 1 114240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_206_421
timestamp 1644511149
transform 1 0 39836 0 1 114240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_206_433
timestamp 1644511149
transform 1 0 40940 0 1 114240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_206_445
timestamp 1644511149
transform 1 0 42044 0 1 114240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_206_457
timestamp 1644511149
transform 1 0 43148 0 1 114240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_206_469
timestamp 1644511149
transform 1 0 44252 0 1 114240
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_206_475
timestamp 1644511149
transform 1 0 44804 0 1 114240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_206_477
timestamp 1644511149
transform 1 0 44988 0 1 114240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_206_489
timestamp 1644511149
transform 1 0 46092 0 1 114240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_206_501
timestamp 1644511149
transform 1 0 47196 0 1 114240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_206_513
timestamp 1644511149
transform 1 0 48300 0 1 114240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_206_525
timestamp 1644511149
transform 1 0 49404 0 1 114240
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_206_531
timestamp 1644511149
transform 1 0 49956 0 1 114240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_206_533
timestamp 1644511149
transform 1 0 50140 0 1 114240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_206_545
timestamp 1644511149
transform 1 0 51244 0 1 114240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_206_557
timestamp 1644511149
transform 1 0 52348 0 1 114240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_206_569
timestamp 1644511149
transform 1 0 53452 0 1 114240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_206_581
timestamp 1644511149
transform 1 0 54556 0 1 114240
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_206_587
timestamp 1644511149
transform 1 0 55108 0 1 114240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_206_589
timestamp 1644511149
transform 1 0 55292 0 1 114240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_206_601
timestamp 1644511149
transform 1 0 56396 0 1 114240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_206_613
timestamp 1644511149
transform 1 0 57500 0 1 114240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_206_625
timestamp 1644511149
transform 1 0 58604 0 1 114240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_206_637
timestamp 1644511149
transform 1 0 59708 0 1 114240
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_206_643
timestamp 1644511149
transform 1 0 60260 0 1 114240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_206_645
timestamp 1644511149
transform 1 0 60444 0 1 114240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_206_657
timestamp 1644511149
transform 1 0 61548 0 1 114240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_206_669
timestamp 1644511149
transform 1 0 62652 0 1 114240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_206_681
timestamp 1644511149
transform 1 0 63756 0 1 114240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_206_693
timestamp 1644511149
transform 1 0 64860 0 1 114240
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_206_699
timestamp 1644511149
transform 1 0 65412 0 1 114240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_206_701
timestamp 1644511149
transform 1 0 65596 0 1 114240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_206_713
timestamp 1644511149
transform 1 0 66700 0 1 114240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_206_725
timestamp 1644511149
transform 1 0 67804 0 1 114240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_206_737
timestamp 1644511149
transform 1 0 68908 0 1 114240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_206_749
timestamp 1644511149
transform 1 0 70012 0 1 114240
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_206_755
timestamp 1644511149
transform 1 0 70564 0 1 114240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_206_757
timestamp 1644511149
transform 1 0 70748 0 1 114240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_206_769
timestamp 1644511149
transform 1 0 71852 0 1 114240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_206_781
timestamp 1644511149
transform 1 0 72956 0 1 114240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_206_793
timestamp 1644511149
transform 1 0 74060 0 1 114240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_206_805
timestamp 1644511149
transform 1 0 75164 0 1 114240
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_206_811
timestamp 1644511149
transform 1 0 75716 0 1 114240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_206_813
timestamp 1644511149
transform 1 0 75900 0 1 114240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_206_825
timestamp 1644511149
transform 1 0 77004 0 1 114240
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_206_833
timestamp 1644511149
transform 1 0 77740 0 1 114240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_206_838
timestamp 1644511149
transform 1 0 78200 0 1 114240
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_207_3
timestamp 1644511149
transform 1 0 1380 0 -1 115328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_207_15
timestamp 1644511149
transform 1 0 2484 0 -1 115328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_207_27
timestamp 1644511149
transform 1 0 3588 0 -1 115328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_207_39
timestamp 1644511149
transform 1 0 4692 0 -1 115328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_207_51
timestamp 1644511149
transform 1 0 5796 0 -1 115328
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_207_55
timestamp 1644511149
transform 1 0 6164 0 -1 115328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_207_57
timestamp 1644511149
transform 1 0 6348 0 -1 115328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_207_69
timestamp 1644511149
transform 1 0 7452 0 -1 115328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_207_81
timestamp 1644511149
transform 1 0 8556 0 -1 115328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_207_93
timestamp 1644511149
transform 1 0 9660 0 -1 115328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_207_105
timestamp 1644511149
transform 1 0 10764 0 -1 115328
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_207_111
timestamp 1644511149
transform 1 0 11316 0 -1 115328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_207_113
timestamp 1644511149
transform 1 0 11500 0 -1 115328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_207_125
timestamp 1644511149
transform 1 0 12604 0 -1 115328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_207_137
timestamp 1644511149
transform 1 0 13708 0 -1 115328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_207_149
timestamp 1644511149
transform 1 0 14812 0 -1 115328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_207_161
timestamp 1644511149
transform 1 0 15916 0 -1 115328
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_207_167
timestamp 1644511149
transform 1 0 16468 0 -1 115328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_207_169
timestamp 1644511149
transform 1 0 16652 0 -1 115328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_207_181
timestamp 1644511149
transform 1 0 17756 0 -1 115328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_207_193
timestamp 1644511149
transform 1 0 18860 0 -1 115328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_207_205
timestamp 1644511149
transform 1 0 19964 0 -1 115328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_207_217
timestamp 1644511149
transform 1 0 21068 0 -1 115328
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_207_223
timestamp 1644511149
transform 1 0 21620 0 -1 115328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_207_225
timestamp 1644511149
transform 1 0 21804 0 -1 115328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_207_237
timestamp 1644511149
transform 1 0 22908 0 -1 115328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_207_249
timestamp 1644511149
transform 1 0 24012 0 -1 115328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_207_261
timestamp 1644511149
transform 1 0 25116 0 -1 115328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_207_273
timestamp 1644511149
transform 1 0 26220 0 -1 115328
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_207_279
timestamp 1644511149
transform 1 0 26772 0 -1 115328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_207_281
timestamp 1644511149
transform 1 0 26956 0 -1 115328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_207_293
timestamp 1644511149
transform 1 0 28060 0 -1 115328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_207_305
timestamp 1644511149
transform 1 0 29164 0 -1 115328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_207_317
timestamp 1644511149
transform 1 0 30268 0 -1 115328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_207_329
timestamp 1644511149
transform 1 0 31372 0 -1 115328
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_207_335
timestamp 1644511149
transform 1 0 31924 0 -1 115328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_207_337
timestamp 1644511149
transform 1 0 32108 0 -1 115328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_207_349
timestamp 1644511149
transform 1 0 33212 0 -1 115328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_207_361
timestamp 1644511149
transform 1 0 34316 0 -1 115328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_207_373
timestamp 1644511149
transform 1 0 35420 0 -1 115328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_207_385
timestamp 1644511149
transform 1 0 36524 0 -1 115328
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_207_391
timestamp 1644511149
transform 1 0 37076 0 -1 115328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_207_393
timestamp 1644511149
transform 1 0 37260 0 -1 115328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_207_405
timestamp 1644511149
transform 1 0 38364 0 -1 115328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_207_417
timestamp 1644511149
transform 1 0 39468 0 -1 115328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_207_429
timestamp 1644511149
transform 1 0 40572 0 -1 115328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_207_441
timestamp 1644511149
transform 1 0 41676 0 -1 115328
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_207_447
timestamp 1644511149
transform 1 0 42228 0 -1 115328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_207_449
timestamp 1644511149
transform 1 0 42412 0 -1 115328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_207_461
timestamp 1644511149
transform 1 0 43516 0 -1 115328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_207_473
timestamp 1644511149
transform 1 0 44620 0 -1 115328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_207_485
timestamp 1644511149
transform 1 0 45724 0 -1 115328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_207_497
timestamp 1644511149
transform 1 0 46828 0 -1 115328
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_207_503
timestamp 1644511149
transform 1 0 47380 0 -1 115328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_207_505
timestamp 1644511149
transform 1 0 47564 0 -1 115328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_207_517
timestamp 1644511149
transform 1 0 48668 0 -1 115328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_207_529
timestamp 1644511149
transform 1 0 49772 0 -1 115328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_207_541
timestamp 1644511149
transform 1 0 50876 0 -1 115328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_207_553
timestamp 1644511149
transform 1 0 51980 0 -1 115328
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_207_559
timestamp 1644511149
transform 1 0 52532 0 -1 115328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_207_561
timestamp 1644511149
transform 1 0 52716 0 -1 115328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_207_573
timestamp 1644511149
transform 1 0 53820 0 -1 115328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_207_585
timestamp 1644511149
transform 1 0 54924 0 -1 115328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_207_597
timestamp 1644511149
transform 1 0 56028 0 -1 115328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_207_609
timestamp 1644511149
transform 1 0 57132 0 -1 115328
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_207_615
timestamp 1644511149
transform 1 0 57684 0 -1 115328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_207_617
timestamp 1644511149
transform 1 0 57868 0 -1 115328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_207_629
timestamp 1644511149
transform 1 0 58972 0 -1 115328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_207_641
timestamp 1644511149
transform 1 0 60076 0 -1 115328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_207_653
timestamp 1644511149
transform 1 0 61180 0 -1 115328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_207_665
timestamp 1644511149
transform 1 0 62284 0 -1 115328
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_207_671
timestamp 1644511149
transform 1 0 62836 0 -1 115328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_207_673
timestamp 1644511149
transform 1 0 63020 0 -1 115328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_207_685
timestamp 1644511149
transform 1 0 64124 0 -1 115328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_207_697
timestamp 1644511149
transform 1 0 65228 0 -1 115328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_207_709
timestamp 1644511149
transform 1 0 66332 0 -1 115328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_207_721
timestamp 1644511149
transform 1 0 67436 0 -1 115328
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_207_727
timestamp 1644511149
transform 1 0 67988 0 -1 115328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_207_729
timestamp 1644511149
transform 1 0 68172 0 -1 115328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_207_741
timestamp 1644511149
transform 1 0 69276 0 -1 115328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_207_753
timestamp 1644511149
transform 1 0 70380 0 -1 115328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_207_765
timestamp 1644511149
transform 1 0 71484 0 -1 115328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_207_777
timestamp 1644511149
transform 1 0 72588 0 -1 115328
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_207_783
timestamp 1644511149
transform 1 0 73140 0 -1 115328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_207_785
timestamp 1644511149
transform 1 0 73324 0 -1 115328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_207_797
timestamp 1644511149
transform 1 0 74428 0 -1 115328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_207_809
timestamp 1644511149
transform 1 0 75532 0 -1 115328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_207_821
timestamp 1644511149
transform 1 0 76636 0 -1 115328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_207_833
timestamp 1644511149
transform 1 0 77740 0 -1 115328
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_207_839
timestamp 1644511149
transform 1 0 78292 0 -1 115328
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_207_841
timestamp 1644511149
transform 1 0 78476 0 -1 115328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_208_3
timestamp 1644511149
transform 1 0 1380 0 1 115328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_208_15
timestamp 1644511149
transform 1 0 2484 0 1 115328
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_208_27
timestamp 1644511149
transform 1 0 3588 0 1 115328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_208_29
timestamp 1644511149
transform 1 0 3772 0 1 115328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_208_41
timestamp 1644511149
transform 1 0 4876 0 1 115328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_208_53
timestamp 1644511149
transform 1 0 5980 0 1 115328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_208_65
timestamp 1644511149
transform 1 0 7084 0 1 115328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_208_77
timestamp 1644511149
transform 1 0 8188 0 1 115328
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_208_83
timestamp 1644511149
transform 1 0 8740 0 1 115328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_208_85
timestamp 1644511149
transform 1 0 8924 0 1 115328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_208_97
timestamp 1644511149
transform 1 0 10028 0 1 115328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_208_109
timestamp 1644511149
transform 1 0 11132 0 1 115328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_208_121
timestamp 1644511149
transform 1 0 12236 0 1 115328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_208_133
timestamp 1644511149
transform 1 0 13340 0 1 115328
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_208_139
timestamp 1644511149
transform 1 0 13892 0 1 115328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_208_141
timestamp 1644511149
transform 1 0 14076 0 1 115328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_208_153
timestamp 1644511149
transform 1 0 15180 0 1 115328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_208_165
timestamp 1644511149
transform 1 0 16284 0 1 115328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_208_177
timestamp 1644511149
transform 1 0 17388 0 1 115328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_208_189
timestamp 1644511149
transform 1 0 18492 0 1 115328
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_208_195
timestamp 1644511149
transform 1 0 19044 0 1 115328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_208_197
timestamp 1644511149
transform 1 0 19228 0 1 115328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_208_209
timestamp 1644511149
transform 1 0 20332 0 1 115328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_208_221
timestamp 1644511149
transform 1 0 21436 0 1 115328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_208_233
timestamp 1644511149
transform 1 0 22540 0 1 115328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_208_245
timestamp 1644511149
transform 1 0 23644 0 1 115328
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_208_251
timestamp 1644511149
transform 1 0 24196 0 1 115328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_208_253
timestamp 1644511149
transform 1 0 24380 0 1 115328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_208_265
timestamp 1644511149
transform 1 0 25484 0 1 115328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_208_277
timestamp 1644511149
transform 1 0 26588 0 1 115328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_208_289
timestamp 1644511149
transform 1 0 27692 0 1 115328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_208_301
timestamp 1644511149
transform 1 0 28796 0 1 115328
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_208_307
timestamp 1644511149
transform 1 0 29348 0 1 115328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_208_309
timestamp 1644511149
transform 1 0 29532 0 1 115328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_208_321
timestamp 1644511149
transform 1 0 30636 0 1 115328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_208_333
timestamp 1644511149
transform 1 0 31740 0 1 115328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_208_345
timestamp 1644511149
transform 1 0 32844 0 1 115328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_208_357
timestamp 1644511149
transform 1 0 33948 0 1 115328
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_208_363
timestamp 1644511149
transform 1 0 34500 0 1 115328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_208_365
timestamp 1644511149
transform 1 0 34684 0 1 115328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_208_377
timestamp 1644511149
transform 1 0 35788 0 1 115328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_208_389
timestamp 1644511149
transform 1 0 36892 0 1 115328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_208_401
timestamp 1644511149
transform 1 0 37996 0 1 115328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_208_413
timestamp 1644511149
transform 1 0 39100 0 1 115328
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_208_419
timestamp 1644511149
transform 1 0 39652 0 1 115328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_208_421
timestamp 1644511149
transform 1 0 39836 0 1 115328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_208_433
timestamp 1644511149
transform 1 0 40940 0 1 115328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_208_445
timestamp 1644511149
transform 1 0 42044 0 1 115328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_208_457
timestamp 1644511149
transform 1 0 43148 0 1 115328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_208_469
timestamp 1644511149
transform 1 0 44252 0 1 115328
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_208_475
timestamp 1644511149
transform 1 0 44804 0 1 115328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_208_477
timestamp 1644511149
transform 1 0 44988 0 1 115328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_208_489
timestamp 1644511149
transform 1 0 46092 0 1 115328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_208_501
timestamp 1644511149
transform 1 0 47196 0 1 115328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_208_513
timestamp 1644511149
transform 1 0 48300 0 1 115328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_208_525
timestamp 1644511149
transform 1 0 49404 0 1 115328
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_208_531
timestamp 1644511149
transform 1 0 49956 0 1 115328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_208_533
timestamp 1644511149
transform 1 0 50140 0 1 115328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_208_545
timestamp 1644511149
transform 1 0 51244 0 1 115328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_208_557
timestamp 1644511149
transform 1 0 52348 0 1 115328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_208_569
timestamp 1644511149
transform 1 0 53452 0 1 115328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_208_581
timestamp 1644511149
transform 1 0 54556 0 1 115328
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_208_587
timestamp 1644511149
transform 1 0 55108 0 1 115328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_208_589
timestamp 1644511149
transform 1 0 55292 0 1 115328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_208_601
timestamp 1644511149
transform 1 0 56396 0 1 115328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_208_613
timestamp 1644511149
transform 1 0 57500 0 1 115328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_208_625
timestamp 1644511149
transform 1 0 58604 0 1 115328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_208_637
timestamp 1644511149
transform 1 0 59708 0 1 115328
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_208_643
timestamp 1644511149
transform 1 0 60260 0 1 115328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_208_645
timestamp 1644511149
transform 1 0 60444 0 1 115328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_208_657
timestamp 1644511149
transform 1 0 61548 0 1 115328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_208_669
timestamp 1644511149
transform 1 0 62652 0 1 115328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_208_681
timestamp 1644511149
transform 1 0 63756 0 1 115328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_208_693
timestamp 1644511149
transform 1 0 64860 0 1 115328
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_208_699
timestamp 1644511149
transform 1 0 65412 0 1 115328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_208_701
timestamp 1644511149
transform 1 0 65596 0 1 115328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_208_713
timestamp 1644511149
transform 1 0 66700 0 1 115328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_208_725
timestamp 1644511149
transform 1 0 67804 0 1 115328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_208_737
timestamp 1644511149
transform 1 0 68908 0 1 115328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_208_749
timestamp 1644511149
transform 1 0 70012 0 1 115328
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_208_755
timestamp 1644511149
transform 1 0 70564 0 1 115328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_208_757
timestamp 1644511149
transform 1 0 70748 0 1 115328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_208_769
timestamp 1644511149
transform 1 0 71852 0 1 115328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_208_781
timestamp 1644511149
transform 1 0 72956 0 1 115328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_208_793
timestamp 1644511149
transform 1 0 74060 0 1 115328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_208_805
timestamp 1644511149
transform 1 0 75164 0 1 115328
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_208_811
timestamp 1644511149
transform 1 0 75716 0 1 115328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_208_813
timestamp 1644511149
transform 1 0 75900 0 1 115328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_208_825
timestamp 1644511149
transform 1 0 77004 0 1 115328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_208_837
timestamp 1644511149
transform 1 0 78108 0 1 115328
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_208_841
timestamp 1644511149
transform 1 0 78476 0 1 115328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_209_3
timestamp 1644511149
transform 1 0 1380 0 -1 116416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_209_15
timestamp 1644511149
transform 1 0 2484 0 -1 116416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_209_27
timestamp 1644511149
transform 1 0 3588 0 -1 116416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_209_39
timestamp 1644511149
transform 1 0 4692 0 -1 116416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_209_51
timestamp 1644511149
transform 1 0 5796 0 -1 116416
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_209_55
timestamp 1644511149
transform 1 0 6164 0 -1 116416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_209_57
timestamp 1644511149
transform 1 0 6348 0 -1 116416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_209_69
timestamp 1644511149
transform 1 0 7452 0 -1 116416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_209_81
timestamp 1644511149
transform 1 0 8556 0 -1 116416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_209_93
timestamp 1644511149
transform 1 0 9660 0 -1 116416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_209_105
timestamp 1644511149
transform 1 0 10764 0 -1 116416
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_209_111
timestamp 1644511149
transform 1 0 11316 0 -1 116416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_209_113
timestamp 1644511149
transform 1 0 11500 0 -1 116416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_209_125
timestamp 1644511149
transform 1 0 12604 0 -1 116416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_209_137
timestamp 1644511149
transform 1 0 13708 0 -1 116416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_209_149
timestamp 1644511149
transform 1 0 14812 0 -1 116416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_209_161
timestamp 1644511149
transform 1 0 15916 0 -1 116416
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_209_167
timestamp 1644511149
transform 1 0 16468 0 -1 116416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_209_169
timestamp 1644511149
transform 1 0 16652 0 -1 116416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_209_181
timestamp 1644511149
transform 1 0 17756 0 -1 116416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_209_193
timestamp 1644511149
transform 1 0 18860 0 -1 116416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_209_205
timestamp 1644511149
transform 1 0 19964 0 -1 116416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_209_217
timestamp 1644511149
transform 1 0 21068 0 -1 116416
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_209_223
timestamp 1644511149
transform 1 0 21620 0 -1 116416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_209_225
timestamp 1644511149
transform 1 0 21804 0 -1 116416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_209_237
timestamp 1644511149
transform 1 0 22908 0 -1 116416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_209_249
timestamp 1644511149
transform 1 0 24012 0 -1 116416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_209_261
timestamp 1644511149
transform 1 0 25116 0 -1 116416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_209_273
timestamp 1644511149
transform 1 0 26220 0 -1 116416
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_209_279
timestamp 1644511149
transform 1 0 26772 0 -1 116416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_209_281
timestamp 1644511149
transform 1 0 26956 0 -1 116416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_209_293
timestamp 1644511149
transform 1 0 28060 0 -1 116416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_209_305
timestamp 1644511149
transform 1 0 29164 0 -1 116416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_209_317
timestamp 1644511149
transform 1 0 30268 0 -1 116416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_209_329
timestamp 1644511149
transform 1 0 31372 0 -1 116416
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_209_335
timestamp 1644511149
transform 1 0 31924 0 -1 116416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_209_337
timestamp 1644511149
transform 1 0 32108 0 -1 116416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_209_349
timestamp 1644511149
transform 1 0 33212 0 -1 116416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_209_361
timestamp 1644511149
transform 1 0 34316 0 -1 116416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_209_373
timestamp 1644511149
transform 1 0 35420 0 -1 116416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_209_385
timestamp 1644511149
transform 1 0 36524 0 -1 116416
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_209_391
timestamp 1644511149
transform 1 0 37076 0 -1 116416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_209_393
timestamp 1644511149
transform 1 0 37260 0 -1 116416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_209_405
timestamp 1644511149
transform 1 0 38364 0 -1 116416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_209_417
timestamp 1644511149
transform 1 0 39468 0 -1 116416
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_209_425
timestamp 1644511149
transform 1 0 40204 0 -1 116416
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_209_433
timestamp 1644511149
transform 1 0 40940 0 -1 116416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_209_445
timestamp 1644511149
transform 1 0 42044 0 -1 116416
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_209_449
timestamp 1644511149
transform 1 0 42412 0 -1 116416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_209_461
timestamp 1644511149
transform 1 0 43516 0 -1 116416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_209_473
timestamp 1644511149
transform 1 0 44620 0 -1 116416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_209_485
timestamp 1644511149
transform 1 0 45724 0 -1 116416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_209_497
timestamp 1644511149
transform 1 0 46828 0 -1 116416
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_209_503
timestamp 1644511149
transform 1 0 47380 0 -1 116416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_209_505
timestamp 1644511149
transform 1 0 47564 0 -1 116416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_209_517
timestamp 1644511149
transform 1 0 48668 0 -1 116416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_209_529
timestamp 1644511149
transform 1 0 49772 0 -1 116416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_209_541
timestamp 1644511149
transform 1 0 50876 0 -1 116416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_209_553
timestamp 1644511149
transform 1 0 51980 0 -1 116416
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_209_559
timestamp 1644511149
transform 1 0 52532 0 -1 116416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_209_561
timestamp 1644511149
transform 1 0 52716 0 -1 116416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_209_573
timestamp 1644511149
transform 1 0 53820 0 -1 116416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_209_585
timestamp 1644511149
transform 1 0 54924 0 -1 116416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_209_597
timestamp 1644511149
transform 1 0 56028 0 -1 116416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_209_609
timestamp 1644511149
transform 1 0 57132 0 -1 116416
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_209_615
timestamp 1644511149
transform 1 0 57684 0 -1 116416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_209_617
timestamp 1644511149
transform 1 0 57868 0 -1 116416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_209_629
timestamp 1644511149
transform 1 0 58972 0 -1 116416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_209_641
timestamp 1644511149
transform 1 0 60076 0 -1 116416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_209_653
timestamp 1644511149
transform 1 0 61180 0 -1 116416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_209_665
timestamp 1644511149
transform 1 0 62284 0 -1 116416
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_209_671
timestamp 1644511149
transform 1 0 62836 0 -1 116416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_209_673
timestamp 1644511149
transform 1 0 63020 0 -1 116416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_209_685
timestamp 1644511149
transform 1 0 64124 0 -1 116416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_209_697
timestamp 1644511149
transform 1 0 65228 0 -1 116416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_209_709
timestamp 1644511149
transform 1 0 66332 0 -1 116416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_209_721
timestamp 1644511149
transform 1 0 67436 0 -1 116416
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_209_727
timestamp 1644511149
transform 1 0 67988 0 -1 116416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_209_729
timestamp 1644511149
transform 1 0 68172 0 -1 116416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_209_741
timestamp 1644511149
transform 1 0 69276 0 -1 116416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_209_753
timestamp 1644511149
transform 1 0 70380 0 -1 116416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_209_765
timestamp 1644511149
transform 1 0 71484 0 -1 116416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_209_777
timestamp 1644511149
transform 1 0 72588 0 -1 116416
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_209_783
timestamp 1644511149
transform 1 0 73140 0 -1 116416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_209_785
timestamp 1644511149
transform 1 0 73324 0 -1 116416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_209_797
timestamp 1644511149
transform 1 0 74428 0 -1 116416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_209_809
timestamp 1644511149
transform 1 0 75532 0 -1 116416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_209_821
timestamp 1644511149
transform 1 0 76636 0 -1 116416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_209_833
timestamp 1644511149
transform 1 0 77740 0 -1 116416
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_209_839
timestamp 1644511149
transform 1 0 78292 0 -1 116416
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_209_841
timestamp 1644511149
transform 1 0 78476 0 -1 116416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_210_3
timestamp 1644511149
transform 1 0 1380 0 1 116416
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_210_13
timestamp 1644511149
transform 1 0 2300 0 1 116416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_210_25
timestamp 1644511149
transform 1 0 3404 0 1 116416
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_210_29
timestamp 1644511149
transform 1 0 3772 0 1 116416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_210_41
timestamp 1644511149
transform 1 0 4876 0 1 116416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_210_53
timestamp 1644511149
transform 1 0 5980 0 1 116416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_210_65
timestamp 1644511149
transform 1 0 7084 0 1 116416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_210_77
timestamp 1644511149
transform 1 0 8188 0 1 116416
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_210_83
timestamp 1644511149
transform 1 0 8740 0 1 116416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_210_85
timestamp 1644511149
transform 1 0 8924 0 1 116416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_210_97
timestamp 1644511149
transform 1 0 10028 0 1 116416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_210_109
timestamp 1644511149
transform 1 0 11132 0 1 116416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_210_121
timestamp 1644511149
transform 1 0 12236 0 1 116416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_210_133
timestamp 1644511149
transform 1 0 13340 0 1 116416
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_210_139
timestamp 1644511149
transform 1 0 13892 0 1 116416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_210_141
timestamp 1644511149
transform 1 0 14076 0 1 116416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_210_153
timestamp 1644511149
transform 1 0 15180 0 1 116416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_210_165
timestamp 1644511149
transform 1 0 16284 0 1 116416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_210_177
timestamp 1644511149
transform 1 0 17388 0 1 116416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_210_189
timestamp 1644511149
transform 1 0 18492 0 1 116416
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_210_195
timestamp 1644511149
transform 1 0 19044 0 1 116416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_210_197
timestamp 1644511149
transform 1 0 19228 0 1 116416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_210_209
timestamp 1644511149
transform 1 0 20332 0 1 116416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_210_221
timestamp 1644511149
transform 1 0 21436 0 1 116416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_210_233
timestamp 1644511149
transform 1 0 22540 0 1 116416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_210_245
timestamp 1644511149
transform 1 0 23644 0 1 116416
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_210_251
timestamp 1644511149
transform 1 0 24196 0 1 116416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_210_253
timestamp 1644511149
transform 1 0 24380 0 1 116416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_210_265
timestamp 1644511149
transform 1 0 25484 0 1 116416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_210_277
timestamp 1644511149
transform 1 0 26588 0 1 116416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_210_289
timestamp 1644511149
transform 1 0 27692 0 1 116416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_210_301
timestamp 1644511149
transform 1 0 28796 0 1 116416
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_210_307
timestamp 1644511149
transform 1 0 29348 0 1 116416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_210_309
timestamp 1644511149
transform 1 0 29532 0 1 116416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_210_321
timestamp 1644511149
transform 1 0 30636 0 1 116416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_210_333
timestamp 1644511149
transform 1 0 31740 0 1 116416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_210_345
timestamp 1644511149
transform 1 0 32844 0 1 116416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_210_357
timestamp 1644511149
transform 1 0 33948 0 1 116416
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_210_363
timestamp 1644511149
transform 1 0 34500 0 1 116416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_210_365
timestamp 1644511149
transform 1 0 34684 0 1 116416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_210_377
timestamp 1644511149
transform 1 0 35788 0 1 116416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_210_389
timestamp 1644511149
transform 1 0 36892 0 1 116416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_210_401
timestamp 1644511149
transform 1 0 37996 0 1 116416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_210_413
timestamp 1644511149
transform 1 0 39100 0 1 116416
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_210_419
timestamp 1644511149
transform 1 0 39652 0 1 116416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_210_421
timestamp 1644511149
transform 1 0 39836 0 1 116416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_210_433
timestamp 1644511149
transform 1 0 40940 0 1 116416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_210_445
timestamp 1644511149
transform 1 0 42044 0 1 116416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_210_457
timestamp 1644511149
transform 1 0 43148 0 1 116416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_210_469
timestamp 1644511149
transform 1 0 44252 0 1 116416
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_210_475
timestamp 1644511149
transform 1 0 44804 0 1 116416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_210_477
timestamp 1644511149
transform 1 0 44988 0 1 116416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_210_489
timestamp 1644511149
transform 1 0 46092 0 1 116416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_210_501
timestamp 1644511149
transform 1 0 47196 0 1 116416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_210_513
timestamp 1644511149
transform 1 0 48300 0 1 116416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_210_525
timestamp 1644511149
transform 1 0 49404 0 1 116416
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_210_531
timestamp 1644511149
transform 1 0 49956 0 1 116416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_210_533
timestamp 1644511149
transform 1 0 50140 0 1 116416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_210_545
timestamp 1644511149
transform 1 0 51244 0 1 116416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_210_557
timestamp 1644511149
transform 1 0 52348 0 1 116416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_210_569
timestamp 1644511149
transform 1 0 53452 0 1 116416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_210_581
timestamp 1644511149
transform 1 0 54556 0 1 116416
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_210_587
timestamp 1644511149
transform 1 0 55108 0 1 116416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_210_589
timestamp 1644511149
transform 1 0 55292 0 1 116416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_210_601
timestamp 1644511149
transform 1 0 56396 0 1 116416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_210_613
timestamp 1644511149
transform 1 0 57500 0 1 116416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_210_625
timestamp 1644511149
transform 1 0 58604 0 1 116416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_210_637
timestamp 1644511149
transform 1 0 59708 0 1 116416
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_210_643
timestamp 1644511149
transform 1 0 60260 0 1 116416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_210_645
timestamp 1644511149
transform 1 0 60444 0 1 116416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_210_657
timestamp 1644511149
transform 1 0 61548 0 1 116416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_210_669
timestamp 1644511149
transform 1 0 62652 0 1 116416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_210_681
timestamp 1644511149
transform 1 0 63756 0 1 116416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_210_693
timestamp 1644511149
transform 1 0 64860 0 1 116416
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_210_699
timestamp 1644511149
transform 1 0 65412 0 1 116416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_210_701
timestamp 1644511149
transform 1 0 65596 0 1 116416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_210_713
timestamp 1644511149
transform 1 0 66700 0 1 116416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_210_725
timestamp 1644511149
transform 1 0 67804 0 1 116416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_210_737
timestamp 1644511149
transform 1 0 68908 0 1 116416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_210_749
timestamp 1644511149
transform 1 0 70012 0 1 116416
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_210_755
timestamp 1644511149
transform 1 0 70564 0 1 116416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_210_757
timestamp 1644511149
transform 1 0 70748 0 1 116416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_210_769
timestamp 1644511149
transform 1 0 71852 0 1 116416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_210_781
timestamp 1644511149
transform 1 0 72956 0 1 116416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_210_793
timestamp 1644511149
transform 1 0 74060 0 1 116416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_210_805
timestamp 1644511149
transform 1 0 75164 0 1 116416
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_210_811
timestamp 1644511149
transform 1 0 75716 0 1 116416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_210_813
timestamp 1644511149
transform 1 0 75900 0 1 116416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_210_825
timestamp 1644511149
transform 1 0 77004 0 1 116416
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_210_833
timestamp 1644511149
transform 1 0 77740 0 1 116416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_210_838
timestamp 1644511149
transform 1 0 78200 0 1 116416
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_211_3
timestamp 1644511149
transform 1 0 1380 0 -1 117504
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_211_13
timestamp 1644511149
transform 1 0 2300 0 -1 117504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_211_25
timestamp 1644511149
transform 1 0 3404 0 -1 117504
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_211_29
timestamp 1644511149
transform 1 0 3772 0 -1 117504
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_211_37
timestamp 1644511149
transform 1 0 4508 0 -1 117504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_211_49
timestamp 1644511149
transform 1 0 5612 0 -1 117504
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_211_55
timestamp 1644511149
transform 1 0 6164 0 -1 117504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_211_57
timestamp 1644511149
transform 1 0 6348 0 -1 117504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_211_69
timestamp 1644511149
transform 1 0 7452 0 -1 117504
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_211_77
timestamp 1644511149
transform 1 0 8188 0 -1 117504
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_211_83
timestamp 1644511149
transform 1 0 8740 0 -1 117504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_211_85
timestamp 1644511149
transform 1 0 8924 0 -1 117504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_211_97
timestamp 1644511149
transform 1 0 10028 0 -1 117504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_211_109
timestamp 1644511149
transform 1 0 11132 0 -1 117504
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_211_113
timestamp 1644511149
transform 1 0 11500 0 -1 117504
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_211_121
timestamp 1644511149
transform 1 0 12236 0 -1 117504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_211_133
timestamp 1644511149
transform 1 0 13340 0 -1 117504
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_211_139
timestamp 1644511149
transform 1 0 13892 0 -1 117504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_211_141
timestamp 1644511149
transform 1 0 14076 0 -1 117504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_211_153
timestamp 1644511149
transform 1 0 15180 0 -1 117504
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_211_161
timestamp 1644511149
transform 1 0 15916 0 -1 117504
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_211_167
timestamp 1644511149
transform 1 0 16468 0 -1 117504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_211_169
timestamp 1644511149
transform 1 0 16652 0 -1 117504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_211_181
timestamp 1644511149
transform 1 0 17756 0 -1 117504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_211_193
timestamp 1644511149
transform 1 0 18860 0 -1 117504
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_211_197
timestamp 1644511149
transform 1 0 19228 0 -1 117504
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_211_203
timestamp 1644511149
transform 1 0 19780 0 -1 117504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_211_215
timestamp 1644511149
transform 1 0 20884 0 -1 117504
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_211_223
timestamp 1644511149
transform 1 0 21620 0 -1 117504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_211_225
timestamp 1644511149
transform 1 0 21804 0 -1 117504
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_211_233
timestamp 1644511149
transform 1 0 22540 0 -1 117504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_211_238
timestamp 1644511149
transform 1 0 23000 0 -1 117504
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_211_250
timestamp 1644511149
transform 1 0 24104 0 -1 117504
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_211_253
timestamp 1644511149
transform 1 0 24380 0 -1 117504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_211_265
timestamp 1644511149
transform 1 0 25484 0 -1 117504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_211_277
timestamp 1644511149
transform 1 0 26588 0 -1 117504
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_211_284
timestamp 1644511149
transform 1 0 27232 0 -1 117504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_211_296
timestamp 1644511149
transform 1 0 28336 0 -1 117504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_211_309
timestamp 1644511149
transform 1 0 29532 0 -1 117504
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_211_317
timestamp 1644511149
transform 1 0 30268 0 -1 117504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_211_322
timestamp 1644511149
transform 1 0 30728 0 -1 117504
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_211_334
timestamp 1644511149
transform 1 0 31832 0 -1 117504
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_211_337
timestamp 1644511149
transform 1 0 32108 0 -1 117504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_211_349
timestamp 1644511149
transform 1 0 33212 0 -1 117504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_211_361
timestamp 1644511149
transform 1 0 34316 0 -1 117504
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_211_369
timestamp 1644511149
transform 1 0 35052 0 -1 117504
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_211_373
timestamp 1644511149
transform 1 0 35420 0 -1 117504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_211_385
timestamp 1644511149
transform 1 0 36524 0 -1 117504
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_211_391
timestamp 1644511149
transform 1 0 37076 0 -1 117504
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_211_393
timestamp 1644511149
transform 1 0 37260 0 -1 117504
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_211_399
timestamp 1644511149
transform 1 0 37812 0 -1 117504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_211_411
timestamp 1644511149
transform 1 0 38916 0 -1 117504
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_211_419
timestamp 1644511149
transform 1 0 39652 0 -1 117504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_211_421
timestamp 1644511149
transform 1 0 39836 0 -1 117504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_211_433
timestamp 1644511149
transform 1 0 40940 0 -1 117504
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_211_441
timestamp 1644511149
transform 1 0 41676 0 -1 117504
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_211_447
timestamp 1644511149
transform 1 0 42228 0 -1 117504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_211_449
timestamp 1644511149
transform 1 0 42412 0 -1 117504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_211_461
timestamp 1644511149
transform 1 0 43516 0 -1 117504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_211_473
timestamp 1644511149
transform 1 0 44620 0 -1 117504
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_211_477
timestamp 1644511149
transform 1 0 44988 0 -1 117504
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_211_483
timestamp 1644511149
transform 1 0 45540 0 -1 117504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_211_495
timestamp 1644511149
transform 1 0 46644 0 -1 117504
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_211_503
timestamp 1644511149
transform 1 0 47380 0 -1 117504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_211_505
timestamp 1644511149
transform 1 0 47564 0 -1 117504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_211_517
timestamp 1644511149
transform 1 0 48668 0 -1 117504
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_211_524
timestamp 1644511149
transform 1 0 49312 0 -1 117504
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_211_533
timestamp 1644511149
transform 1 0 50140 0 -1 117504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_211_545
timestamp 1644511149
transform 1 0 51244 0 -1 117504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_211_557
timestamp 1644511149
transform 1 0 52348 0 -1 117504
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_211_565
timestamp 1644511149
transform 1 0 53084 0 -1 117504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_211_577
timestamp 1644511149
transform 1 0 54188 0 -1 117504
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_211_585
timestamp 1644511149
transform 1 0 54924 0 -1 117504
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_211_589
timestamp 1644511149
transform 1 0 55292 0 -1 117504
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_211_597
timestamp 1644511149
transform 1 0 56028 0 -1 117504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_211_604
timestamp 1644511149
transform 1 0 56672 0 -1 117504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_211_617
timestamp 1644511149
transform 1 0 57868 0 -1 117504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_211_629
timestamp 1644511149
transform 1 0 58972 0 -1 117504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_211_641
timestamp 1644511149
transform 1 0 60076 0 -1 117504
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_211_648
timestamp 1644511149
transform 1 0 60720 0 -1 117504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_211_660
timestamp 1644511149
transform 1 0 61824 0 -1 117504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_211_673
timestamp 1644511149
transform 1 0 63020 0 -1 117504
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_211_681
timestamp 1644511149
transform 1 0 63756 0 -1 117504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_211_686
timestamp 1644511149
transform 1 0 64216 0 -1 117504
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_211_698
timestamp 1644511149
transform 1 0 65320 0 -1 117504
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_211_701
timestamp 1644511149
transform 1 0 65596 0 -1 117504
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_211_715
timestamp 1644511149
transform 1 0 66884 0 -1 117504
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_211_721
timestamp 1644511149
transform 1 0 67436 0 -1 117504
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_211_727
timestamp 1644511149
transform 1 0 67988 0 -1 117504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_211_729
timestamp 1644511149
transform 1 0 68172 0 -1 117504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_211_741
timestamp 1644511149
transform 1 0 69276 0 -1 117504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_211_753
timestamp 1644511149
transform 1 0 70380 0 -1 117504
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_211_757
timestamp 1644511149
transform 1 0 70748 0 -1 117504
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_211_767
timestamp 1644511149
transform 1 0 71668 0 -1 117504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_211_779
timestamp 1644511149
transform 1 0 72772 0 -1 117504
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_211_783
timestamp 1644511149
transform 1 0 73140 0 -1 117504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_211_785
timestamp 1644511149
transform 1 0 73324 0 -1 117504
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_211_799
timestamp 1644511149
transform 1 0 74612 0 -1 117504
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_211_805
timestamp 1644511149
transform 1 0 75164 0 -1 117504
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_211_811
timestamp 1644511149
transform 1 0 75716 0 -1 117504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_211_813
timestamp 1644511149
transform 1 0 75900 0 -1 117504
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_211_825
timestamp 1644511149
transform 1 0 77004 0 -1 117504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_211_836
timestamp 1644511149
transform 1 0 78016 0 -1 117504
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_211_841
timestamp 1644511149
transform 1 0 78476 0 -1 117504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1644511149
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1644511149
transform -1 0 78844 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1644511149
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1644511149
transform -1 0 78844 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1644511149
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1644511149
transform -1 0 78844 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1644511149
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1644511149
transform -1 0 78844 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1644511149
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1644511149
transform -1 0 78844 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1644511149
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1644511149
transform -1 0 78844 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1644511149
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1644511149
transform -1 0 78844 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1644511149
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1644511149
transform -1 0 78844 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1644511149
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1644511149
transform -1 0 78844 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1644511149
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1644511149
transform -1 0 78844 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1644511149
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1644511149
transform -1 0 78844 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1644511149
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1644511149
transform -1 0 78844 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1644511149
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1644511149
transform -1 0 78844 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1644511149
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1644511149
transform -1 0 78844 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1644511149
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1644511149
transform -1 0 78844 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1644511149
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1644511149
transform -1 0 78844 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1644511149
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1644511149
transform -1 0 78844 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1644511149
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1644511149
transform -1 0 78844 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1644511149
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1644511149
transform -1 0 78844 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1644511149
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1644511149
transform -1 0 78844 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1644511149
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1644511149
transform -1 0 78844 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1644511149
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1644511149
transform -1 0 78844 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1644511149
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1644511149
transform -1 0 78844 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1644511149
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1644511149
transform -1 0 78844 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1644511149
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1644511149
transform -1 0 78844 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1644511149
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1644511149
transform -1 0 78844 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1644511149
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1644511149
transform -1 0 78844 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1644511149
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1644511149
transform -1 0 78844 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1644511149
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1644511149
transform -1 0 78844 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1644511149
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1644511149
transform -1 0 78844 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1644511149
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1644511149
transform -1 0 78844 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1644511149
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1644511149
transform -1 0 78844 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1644511149
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1644511149
transform -1 0 78844 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1644511149
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1644511149
transform -1 0 78844 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1644511149
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1644511149
transform -1 0 78844 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1644511149
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1644511149
transform -1 0 78844 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1644511149
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1644511149
transform -1 0 78844 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1644511149
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1644511149
transform -1 0 78844 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1644511149
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1644511149
transform -1 0 78844 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1644511149
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1644511149
transform -1 0 78844 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1644511149
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1644511149
transform -1 0 78844 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1644511149
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1644511149
transform -1 0 78844 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1644511149
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1644511149
transform -1 0 78844 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1644511149
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1644511149
transform -1 0 78844 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1644511149
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1644511149
transform -1 0 78844 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1644511149
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1644511149
transform -1 0 78844 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1644511149
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1644511149
transform -1 0 78844 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1644511149
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1644511149
transform -1 0 78844 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1644511149
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1644511149
transform -1 0 78844 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1644511149
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1644511149
transform -1 0 78844 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1644511149
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1644511149
transform -1 0 78844 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1644511149
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1644511149
transform -1 0 78844 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1644511149
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1644511149
transform -1 0 78844 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1644511149
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1644511149
transform -1 0 78844 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1644511149
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1644511149
transform -1 0 78844 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1644511149
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1644511149
transform -1 0 78844 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1644511149
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1644511149
transform -1 0 78844 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1644511149
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1644511149
transform -1 0 78844 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1644511149
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1644511149
transform -1 0 78844 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1644511149
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1644511149
transform -1 0 78844 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1644511149
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1644511149
transform -1 0 78844 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1644511149
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1644511149
transform -1 0 78844 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1644511149
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1644511149
transform -1 0 78844 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1644511149
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1644511149
transform -1 0 78844 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1644511149
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1644511149
transform -1 0 78844 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1644511149
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1644511149
transform -1 0 78844 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1644511149
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1644511149
transform -1 0 78844 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 1644511149
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 1644511149
transform -1 0 78844 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_136
timestamp 1644511149
transform 1 0 1104 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_137
timestamp 1644511149
transform -1 0 78844 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_138
timestamp 1644511149
transform 1 0 1104 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_139
timestamp 1644511149
transform -1 0 78844 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_140
timestamp 1644511149
transform 1 0 1104 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_141
timestamp 1644511149
transform -1 0 78844 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_142
timestamp 1644511149
transform 1 0 1104 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_143
timestamp 1644511149
transform -1 0 78844 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_144
timestamp 1644511149
transform 1 0 1104 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_145
timestamp 1644511149
transform -1 0 78844 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_146
timestamp 1644511149
transform 1 0 1104 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_147
timestamp 1644511149
transform -1 0 78844 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_148
timestamp 1644511149
transform 1 0 1104 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_149
timestamp 1644511149
transform -1 0 78844 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_150
timestamp 1644511149
transform 1 0 1104 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_151
timestamp 1644511149
transform -1 0 78844 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_152
timestamp 1644511149
transform 1 0 1104 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_153
timestamp 1644511149
transform -1 0 78844 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_154
timestamp 1644511149
transform 1 0 1104 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_155
timestamp 1644511149
transform -1 0 78844 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_156
timestamp 1644511149
transform 1 0 1104 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_157
timestamp 1644511149
transform -1 0 78844 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_158
timestamp 1644511149
transform 1 0 1104 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_159
timestamp 1644511149
transform -1 0 78844 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_160
timestamp 1644511149
transform 1 0 1104 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_161
timestamp 1644511149
transform -1 0 78844 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_162
timestamp 1644511149
transform 1 0 1104 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_163
timestamp 1644511149
transform -1 0 78844 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_164
timestamp 1644511149
transform 1 0 1104 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_165
timestamp 1644511149
transform -1 0 78844 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_166
timestamp 1644511149
transform 1 0 1104 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_167
timestamp 1644511149
transform -1 0 78844 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_168
timestamp 1644511149
transform 1 0 1104 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_169
timestamp 1644511149
transform -1 0 78844 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_170
timestamp 1644511149
transform 1 0 1104 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_171
timestamp 1644511149
transform -1 0 78844 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_172
timestamp 1644511149
transform 1 0 1104 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_173
timestamp 1644511149
transform -1 0 78844 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_174
timestamp 1644511149
transform 1 0 1104 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_175
timestamp 1644511149
transform -1 0 78844 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_176
timestamp 1644511149
transform 1 0 1104 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_177
timestamp 1644511149
transform -1 0 78844 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_178
timestamp 1644511149
transform 1 0 1104 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_179
timestamp 1644511149
transform -1 0 78844 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_180
timestamp 1644511149
transform 1 0 1104 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_181
timestamp 1644511149
transform -1 0 78844 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_182
timestamp 1644511149
transform 1 0 1104 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_183
timestamp 1644511149
transform -1 0 78844 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_184
timestamp 1644511149
transform 1 0 1104 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_185
timestamp 1644511149
transform -1 0 78844 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_186
timestamp 1644511149
transform 1 0 1104 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_187
timestamp 1644511149
transform -1 0 78844 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_188
timestamp 1644511149
transform 1 0 1104 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_189
timestamp 1644511149
transform -1 0 78844 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_190
timestamp 1644511149
transform 1 0 1104 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_191
timestamp 1644511149
transform -1 0 78844 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_192
timestamp 1644511149
transform 1 0 1104 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_193
timestamp 1644511149
transform -1 0 78844 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_194
timestamp 1644511149
transform 1 0 1104 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_195
timestamp 1644511149
transform -1 0 78844 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_196
timestamp 1644511149
transform 1 0 1104 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_197
timestamp 1644511149
transform -1 0 78844 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_198
timestamp 1644511149
transform 1 0 1104 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_199
timestamp 1644511149
transform -1 0 78844 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_200
timestamp 1644511149
transform 1 0 1104 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_201
timestamp 1644511149
transform -1 0 78844 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_202
timestamp 1644511149
transform 1 0 1104 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_203
timestamp 1644511149
transform -1 0 78844 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_204
timestamp 1644511149
transform 1 0 1104 0 1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_205
timestamp 1644511149
transform -1 0 78844 0 1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_206
timestamp 1644511149
transform 1 0 1104 0 -1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_207
timestamp 1644511149
transform -1 0 78844 0 -1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_208
timestamp 1644511149
transform 1 0 1104 0 1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_209
timestamp 1644511149
transform -1 0 78844 0 1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_210
timestamp 1644511149
transform 1 0 1104 0 -1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_211
timestamp 1644511149
transform -1 0 78844 0 -1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_212
timestamp 1644511149
transform 1 0 1104 0 1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_213
timestamp 1644511149
transform -1 0 78844 0 1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_214
timestamp 1644511149
transform 1 0 1104 0 -1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_215
timestamp 1644511149
transform -1 0 78844 0 -1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_216
timestamp 1644511149
transform 1 0 1104 0 1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_217
timestamp 1644511149
transform -1 0 78844 0 1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_218
timestamp 1644511149
transform 1 0 1104 0 -1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_219
timestamp 1644511149
transform -1 0 78844 0 -1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_220
timestamp 1644511149
transform 1 0 1104 0 1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_221
timestamp 1644511149
transform -1 0 78844 0 1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_222
timestamp 1644511149
transform 1 0 1104 0 -1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_223
timestamp 1644511149
transform -1 0 78844 0 -1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_224
timestamp 1644511149
transform 1 0 1104 0 1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_225
timestamp 1644511149
transform -1 0 78844 0 1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_226
timestamp 1644511149
transform 1 0 1104 0 -1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_227
timestamp 1644511149
transform -1 0 78844 0 -1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_228
timestamp 1644511149
transform 1 0 1104 0 1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_229
timestamp 1644511149
transform -1 0 78844 0 1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_230
timestamp 1644511149
transform 1 0 1104 0 -1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_231
timestamp 1644511149
transform -1 0 78844 0 -1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_232
timestamp 1644511149
transform 1 0 1104 0 1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_233
timestamp 1644511149
transform -1 0 78844 0 1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_234
timestamp 1644511149
transform 1 0 1104 0 -1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_235
timestamp 1644511149
transform -1 0 78844 0 -1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_236
timestamp 1644511149
transform 1 0 1104 0 1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_237
timestamp 1644511149
transform -1 0 78844 0 1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_238
timestamp 1644511149
transform 1 0 1104 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_239
timestamp 1644511149
transform -1 0 78844 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_240
timestamp 1644511149
transform 1 0 1104 0 1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_241
timestamp 1644511149
transform -1 0 78844 0 1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_242
timestamp 1644511149
transform 1 0 1104 0 -1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_243
timestamp 1644511149
transform -1 0 78844 0 -1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_244
timestamp 1644511149
transform 1 0 1104 0 1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_245
timestamp 1644511149
transform -1 0 78844 0 1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_246
timestamp 1644511149
transform 1 0 1104 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_247
timestamp 1644511149
transform -1 0 78844 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_248
timestamp 1644511149
transform 1 0 1104 0 1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_249
timestamp 1644511149
transform -1 0 78844 0 1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_250
timestamp 1644511149
transform 1 0 1104 0 -1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_251
timestamp 1644511149
transform -1 0 78844 0 -1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_252
timestamp 1644511149
transform 1 0 1104 0 1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_253
timestamp 1644511149
transform -1 0 78844 0 1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_254
timestamp 1644511149
transform 1 0 1104 0 -1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_255
timestamp 1644511149
transform -1 0 78844 0 -1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_256
timestamp 1644511149
transform 1 0 1104 0 1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_257
timestamp 1644511149
transform -1 0 78844 0 1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_258
timestamp 1644511149
transform 1 0 1104 0 -1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_259
timestamp 1644511149
transform -1 0 78844 0 -1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_260
timestamp 1644511149
transform 1 0 1104 0 1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_261
timestamp 1644511149
transform -1 0 78844 0 1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_262
timestamp 1644511149
transform 1 0 1104 0 -1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_263
timestamp 1644511149
transform -1 0 78844 0 -1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_264
timestamp 1644511149
transform 1 0 1104 0 1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_265
timestamp 1644511149
transform -1 0 78844 0 1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_266
timestamp 1644511149
transform 1 0 1104 0 -1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_267
timestamp 1644511149
transform -1 0 78844 0 -1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_268
timestamp 1644511149
transform 1 0 1104 0 1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_269
timestamp 1644511149
transform -1 0 78844 0 1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_270
timestamp 1644511149
transform 1 0 1104 0 -1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_271
timestamp 1644511149
transform -1 0 78844 0 -1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_272
timestamp 1644511149
transform 1 0 1104 0 1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_273
timestamp 1644511149
transform -1 0 78844 0 1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_274
timestamp 1644511149
transform 1 0 1104 0 -1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_275
timestamp 1644511149
transform -1 0 78844 0 -1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_276
timestamp 1644511149
transform 1 0 1104 0 1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_277
timestamp 1644511149
transform -1 0 78844 0 1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_278
timestamp 1644511149
transform 1 0 1104 0 -1 78336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_279
timestamp 1644511149
transform -1 0 78844 0 -1 78336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_280
timestamp 1644511149
transform 1 0 1104 0 1 78336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_281
timestamp 1644511149
transform -1 0 78844 0 1 78336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_282
timestamp 1644511149
transform 1 0 1104 0 -1 79424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_283
timestamp 1644511149
transform -1 0 78844 0 -1 79424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_284
timestamp 1644511149
transform 1 0 1104 0 1 79424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_285
timestamp 1644511149
transform -1 0 78844 0 1 79424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_286
timestamp 1644511149
transform 1 0 1104 0 -1 80512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_287
timestamp 1644511149
transform -1 0 78844 0 -1 80512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_288
timestamp 1644511149
transform 1 0 1104 0 1 80512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_289
timestamp 1644511149
transform -1 0 78844 0 1 80512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_290
timestamp 1644511149
transform 1 0 1104 0 -1 81600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_291
timestamp 1644511149
transform -1 0 78844 0 -1 81600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_292
timestamp 1644511149
transform 1 0 1104 0 1 81600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_293
timestamp 1644511149
transform -1 0 78844 0 1 81600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_294
timestamp 1644511149
transform 1 0 1104 0 -1 82688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_295
timestamp 1644511149
transform -1 0 78844 0 -1 82688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_296
timestamp 1644511149
transform 1 0 1104 0 1 82688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_297
timestamp 1644511149
transform -1 0 78844 0 1 82688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_298
timestamp 1644511149
transform 1 0 1104 0 -1 83776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_299
timestamp 1644511149
transform -1 0 78844 0 -1 83776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_300
timestamp 1644511149
transform 1 0 1104 0 1 83776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_301
timestamp 1644511149
transform -1 0 78844 0 1 83776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_302
timestamp 1644511149
transform 1 0 1104 0 -1 84864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_303
timestamp 1644511149
transform -1 0 78844 0 -1 84864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_304
timestamp 1644511149
transform 1 0 1104 0 1 84864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_305
timestamp 1644511149
transform -1 0 78844 0 1 84864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_306
timestamp 1644511149
transform 1 0 1104 0 -1 85952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_307
timestamp 1644511149
transform -1 0 78844 0 -1 85952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_308
timestamp 1644511149
transform 1 0 1104 0 1 85952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_309
timestamp 1644511149
transform -1 0 78844 0 1 85952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_310
timestamp 1644511149
transform 1 0 1104 0 -1 87040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_311
timestamp 1644511149
transform -1 0 78844 0 -1 87040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_312
timestamp 1644511149
transform 1 0 1104 0 1 87040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_313
timestamp 1644511149
transform -1 0 78844 0 1 87040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_314
timestamp 1644511149
transform 1 0 1104 0 -1 88128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_315
timestamp 1644511149
transform -1 0 78844 0 -1 88128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_316
timestamp 1644511149
transform 1 0 1104 0 1 88128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_317
timestamp 1644511149
transform -1 0 78844 0 1 88128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_318
timestamp 1644511149
transform 1 0 1104 0 -1 89216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_319
timestamp 1644511149
transform -1 0 78844 0 -1 89216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_320
timestamp 1644511149
transform 1 0 1104 0 1 89216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_321
timestamp 1644511149
transform -1 0 78844 0 1 89216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_322
timestamp 1644511149
transform 1 0 1104 0 -1 90304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_323
timestamp 1644511149
transform -1 0 78844 0 -1 90304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_324
timestamp 1644511149
transform 1 0 1104 0 1 90304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_325
timestamp 1644511149
transform -1 0 78844 0 1 90304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_326
timestamp 1644511149
transform 1 0 1104 0 -1 91392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_327
timestamp 1644511149
transform -1 0 78844 0 -1 91392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_328
timestamp 1644511149
transform 1 0 1104 0 1 91392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_329
timestamp 1644511149
transform -1 0 78844 0 1 91392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_330
timestamp 1644511149
transform 1 0 1104 0 -1 92480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_331
timestamp 1644511149
transform -1 0 78844 0 -1 92480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_332
timestamp 1644511149
transform 1 0 1104 0 1 92480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_333
timestamp 1644511149
transform -1 0 78844 0 1 92480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_334
timestamp 1644511149
transform 1 0 1104 0 -1 93568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_335
timestamp 1644511149
transform -1 0 78844 0 -1 93568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_336
timestamp 1644511149
transform 1 0 1104 0 1 93568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_337
timestamp 1644511149
transform -1 0 78844 0 1 93568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_338
timestamp 1644511149
transform 1 0 1104 0 -1 94656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_339
timestamp 1644511149
transform -1 0 78844 0 -1 94656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_340
timestamp 1644511149
transform 1 0 1104 0 1 94656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_341
timestamp 1644511149
transform -1 0 78844 0 1 94656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_342
timestamp 1644511149
transform 1 0 1104 0 -1 95744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_343
timestamp 1644511149
transform -1 0 78844 0 -1 95744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_344
timestamp 1644511149
transform 1 0 1104 0 1 95744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_345
timestamp 1644511149
transform -1 0 78844 0 1 95744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_346
timestamp 1644511149
transform 1 0 1104 0 -1 96832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_347
timestamp 1644511149
transform -1 0 78844 0 -1 96832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_348
timestamp 1644511149
transform 1 0 1104 0 1 96832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_349
timestamp 1644511149
transform -1 0 78844 0 1 96832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_350
timestamp 1644511149
transform 1 0 1104 0 -1 97920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_351
timestamp 1644511149
transform -1 0 78844 0 -1 97920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_352
timestamp 1644511149
transform 1 0 1104 0 1 97920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_353
timestamp 1644511149
transform -1 0 78844 0 1 97920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_354
timestamp 1644511149
transform 1 0 1104 0 -1 99008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_355
timestamp 1644511149
transform -1 0 78844 0 -1 99008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_356
timestamp 1644511149
transform 1 0 1104 0 1 99008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_357
timestamp 1644511149
transform -1 0 78844 0 1 99008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_358
timestamp 1644511149
transform 1 0 1104 0 -1 100096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_359
timestamp 1644511149
transform -1 0 78844 0 -1 100096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_360
timestamp 1644511149
transform 1 0 1104 0 1 100096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_361
timestamp 1644511149
transform -1 0 78844 0 1 100096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_362
timestamp 1644511149
transform 1 0 1104 0 -1 101184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_363
timestamp 1644511149
transform -1 0 78844 0 -1 101184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_364
timestamp 1644511149
transform 1 0 1104 0 1 101184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_365
timestamp 1644511149
transform -1 0 78844 0 1 101184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_366
timestamp 1644511149
transform 1 0 1104 0 -1 102272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_367
timestamp 1644511149
transform -1 0 78844 0 -1 102272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_368
timestamp 1644511149
transform 1 0 1104 0 1 102272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_369
timestamp 1644511149
transform -1 0 78844 0 1 102272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_370
timestamp 1644511149
transform 1 0 1104 0 -1 103360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_371
timestamp 1644511149
transform -1 0 78844 0 -1 103360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_372
timestamp 1644511149
transform 1 0 1104 0 1 103360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_373
timestamp 1644511149
transform -1 0 78844 0 1 103360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_374
timestamp 1644511149
transform 1 0 1104 0 -1 104448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_375
timestamp 1644511149
transform -1 0 78844 0 -1 104448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_376
timestamp 1644511149
transform 1 0 1104 0 1 104448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_377
timestamp 1644511149
transform -1 0 78844 0 1 104448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_378
timestamp 1644511149
transform 1 0 1104 0 -1 105536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_379
timestamp 1644511149
transform -1 0 78844 0 -1 105536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_380
timestamp 1644511149
transform 1 0 1104 0 1 105536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_381
timestamp 1644511149
transform -1 0 78844 0 1 105536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_382
timestamp 1644511149
transform 1 0 1104 0 -1 106624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_383
timestamp 1644511149
transform -1 0 78844 0 -1 106624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_384
timestamp 1644511149
transform 1 0 1104 0 1 106624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_385
timestamp 1644511149
transform -1 0 78844 0 1 106624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_386
timestamp 1644511149
transform 1 0 1104 0 -1 107712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_387
timestamp 1644511149
transform -1 0 78844 0 -1 107712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_388
timestamp 1644511149
transform 1 0 1104 0 1 107712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_389
timestamp 1644511149
transform -1 0 78844 0 1 107712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_390
timestamp 1644511149
transform 1 0 1104 0 -1 108800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_391
timestamp 1644511149
transform -1 0 78844 0 -1 108800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_392
timestamp 1644511149
transform 1 0 1104 0 1 108800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_393
timestamp 1644511149
transform -1 0 78844 0 1 108800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_394
timestamp 1644511149
transform 1 0 1104 0 -1 109888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_395
timestamp 1644511149
transform -1 0 78844 0 -1 109888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_396
timestamp 1644511149
transform 1 0 1104 0 1 109888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_397
timestamp 1644511149
transform -1 0 78844 0 1 109888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_398
timestamp 1644511149
transform 1 0 1104 0 -1 110976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_399
timestamp 1644511149
transform -1 0 78844 0 -1 110976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_400
timestamp 1644511149
transform 1 0 1104 0 1 110976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_401
timestamp 1644511149
transform -1 0 78844 0 1 110976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_402
timestamp 1644511149
transform 1 0 1104 0 -1 112064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_403
timestamp 1644511149
transform -1 0 78844 0 -1 112064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_404
timestamp 1644511149
transform 1 0 1104 0 1 112064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_405
timestamp 1644511149
transform -1 0 78844 0 1 112064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_406
timestamp 1644511149
transform 1 0 1104 0 -1 113152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_407
timestamp 1644511149
transform -1 0 78844 0 -1 113152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_408
timestamp 1644511149
transform 1 0 1104 0 1 113152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_409
timestamp 1644511149
transform -1 0 78844 0 1 113152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_410
timestamp 1644511149
transform 1 0 1104 0 -1 114240
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_411
timestamp 1644511149
transform -1 0 78844 0 -1 114240
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_412
timestamp 1644511149
transform 1 0 1104 0 1 114240
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_413
timestamp 1644511149
transform -1 0 78844 0 1 114240
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_414
timestamp 1644511149
transform 1 0 1104 0 -1 115328
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_415
timestamp 1644511149
transform -1 0 78844 0 -1 115328
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_416
timestamp 1644511149
transform 1 0 1104 0 1 115328
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_417
timestamp 1644511149
transform -1 0 78844 0 1 115328
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_418
timestamp 1644511149
transform 1 0 1104 0 -1 116416
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_419
timestamp 1644511149
transform -1 0 78844 0 -1 116416
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_420
timestamp 1644511149
transform 1 0 1104 0 1 116416
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_421
timestamp 1644511149
transform -1 0 78844 0 1 116416
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_422
timestamp 1644511149
transform 1 0 1104 0 -1 117504
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_423
timestamp 1644511149
transform -1 0 78844 0 -1 117504
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424 caravel_pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1644511149
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1644511149
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1644511149
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1644511149
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1644511149
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1644511149
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1644511149
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1644511149
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1644511149
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1644511149
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1644511149
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1644511149
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1644511149
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1644511149
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1644511149
transform 1 0 42320 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1644511149
transform 1 0 44896 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1644511149
transform 1 0 47472 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1644511149
transform 1 0 50048 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1644511149
transform 1 0 52624 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1644511149
transform 1 0 55200 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1644511149
transform 1 0 57776 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1644511149
transform 1 0 60352 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1644511149
transform 1 0 62928 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1644511149
transform 1 0 65504 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1644511149
transform 1 0 68080 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1644511149
transform 1 0 70656 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1644511149
transform 1 0 73232 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1644511149
transform 1 0 75808 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1644511149
transform 1 0 78384 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1644511149
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1644511149
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1644511149
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1644511149
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1644511149
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1644511149
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1644511149
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1644511149
transform 1 0 42320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1644511149
transform 1 0 47472 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1644511149
transform 1 0 52624 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1644511149
transform 1 0 57776 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1644511149
transform 1 0 62928 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1644511149
transform 1 0 68080 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1644511149
transform 1 0 73232 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1644511149
transform 1 0 78384 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1644511149
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1644511149
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1644511149
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1644511149
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1644511149
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1644511149
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1644511149
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1644511149
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1644511149
transform 1 0 44896 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1644511149
transform 1 0 50048 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1644511149
transform 1 0 55200 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1644511149
transform 1 0 60352 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1644511149
transform 1 0 65504 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1644511149
transform 1 0 70656 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1644511149
transform 1 0 75808 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1644511149
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1644511149
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1644511149
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1644511149
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1644511149
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1644511149
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1644511149
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1644511149
transform 1 0 42320 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1644511149
transform 1 0 47472 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1644511149
transform 1 0 52624 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1644511149
transform 1 0 57776 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1644511149
transform 1 0 62928 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1644511149
transform 1 0 68080 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1644511149
transform 1 0 73232 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1644511149
transform 1 0 78384 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1644511149
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1644511149
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1644511149
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1644511149
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1644511149
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1644511149
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1644511149
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1644511149
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1644511149
transform 1 0 44896 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1644511149
transform 1 0 50048 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1644511149
transform 1 0 55200 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1644511149
transform 1 0 60352 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1644511149
transform 1 0 65504 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1644511149
transform 1 0 70656 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1644511149
transform 1 0 75808 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1644511149
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1644511149
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1644511149
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1644511149
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1644511149
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1644511149
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1644511149
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1644511149
transform 1 0 42320 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1644511149
transform 1 0 47472 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1644511149
transform 1 0 52624 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1644511149
transform 1 0 57776 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1644511149
transform 1 0 62928 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1644511149
transform 1 0 68080 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1644511149
transform 1 0 73232 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1644511149
transform 1 0 78384 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1644511149
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1644511149
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1644511149
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1644511149
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1644511149
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1644511149
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1644511149
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1644511149
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1644511149
transform 1 0 44896 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1644511149
transform 1 0 50048 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1644511149
transform 1 0 55200 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1644511149
transform 1 0 60352 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1644511149
transform 1 0 65504 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1644511149
transform 1 0 70656 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1644511149
transform 1 0 75808 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1644511149
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1644511149
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1644511149
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1644511149
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1644511149
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1644511149
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1644511149
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1644511149
transform 1 0 42320 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1644511149
transform 1 0 47472 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1644511149
transform 1 0 52624 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1644511149
transform 1 0 57776 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1644511149
transform 1 0 62928 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1644511149
transform 1 0 68080 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1644511149
transform 1 0 73232 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1644511149
transform 1 0 78384 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1644511149
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1644511149
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1644511149
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1644511149
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1644511149
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1644511149
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1644511149
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1644511149
transform 1 0 39744 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1644511149
transform 1 0 44896 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1644511149
transform 1 0 50048 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1644511149
transform 1 0 55200 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1644511149
transform 1 0 60352 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1644511149
transform 1 0 65504 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1644511149
transform 1 0 70656 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1644511149
transform 1 0 75808 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1644511149
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1644511149
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1644511149
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1644511149
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1644511149
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1644511149
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1644511149
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1644511149
transform 1 0 42320 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1644511149
transform 1 0 47472 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1644511149
transform 1 0 52624 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1644511149
transform 1 0 57776 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1644511149
transform 1 0 62928 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1644511149
transform 1 0 68080 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1644511149
transform 1 0 73232 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1644511149
transform 1 0 78384 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1644511149
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1644511149
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1644511149
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1644511149
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1644511149
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1644511149
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1644511149
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1644511149
transform 1 0 39744 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1644511149
transform 1 0 44896 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1644511149
transform 1 0 50048 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_599
timestamp 1644511149
transform 1 0 55200 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_600
timestamp 1644511149
transform 1 0 60352 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_601
timestamp 1644511149
transform 1 0 65504 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_602
timestamp 1644511149
transform 1 0 70656 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_603
timestamp 1644511149
transform 1 0 75808 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_604
timestamp 1644511149
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_605
timestamp 1644511149
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_606
timestamp 1644511149
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_607
timestamp 1644511149
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_608
timestamp 1644511149
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_609
timestamp 1644511149
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_610
timestamp 1644511149
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_611
timestamp 1644511149
transform 1 0 42320 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_612
timestamp 1644511149
transform 1 0 47472 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_613
timestamp 1644511149
transform 1 0 52624 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_614
timestamp 1644511149
transform 1 0 57776 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_615
timestamp 1644511149
transform 1 0 62928 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_616
timestamp 1644511149
transform 1 0 68080 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_617
timestamp 1644511149
transform 1 0 73232 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_618
timestamp 1644511149
transform 1 0 78384 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_619
timestamp 1644511149
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_620
timestamp 1644511149
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_621
timestamp 1644511149
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_622
timestamp 1644511149
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_623
timestamp 1644511149
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_624
timestamp 1644511149
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_625
timestamp 1644511149
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_626
timestamp 1644511149
transform 1 0 39744 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_627
timestamp 1644511149
transform 1 0 44896 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_628
timestamp 1644511149
transform 1 0 50048 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_629
timestamp 1644511149
transform 1 0 55200 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_630
timestamp 1644511149
transform 1 0 60352 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_631
timestamp 1644511149
transform 1 0 65504 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_632
timestamp 1644511149
transform 1 0 70656 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_633
timestamp 1644511149
transform 1 0 75808 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_634
timestamp 1644511149
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_635
timestamp 1644511149
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_636
timestamp 1644511149
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_637
timestamp 1644511149
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_638
timestamp 1644511149
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_639
timestamp 1644511149
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_640
timestamp 1644511149
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_641
timestamp 1644511149
transform 1 0 42320 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_642
timestamp 1644511149
transform 1 0 47472 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_643
timestamp 1644511149
transform 1 0 52624 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_644
timestamp 1644511149
transform 1 0 57776 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_645
timestamp 1644511149
transform 1 0 62928 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_646
timestamp 1644511149
transform 1 0 68080 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_647
timestamp 1644511149
transform 1 0 73232 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_648
timestamp 1644511149
transform 1 0 78384 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_649
timestamp 1644511149
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_650
timestamp 1644511149
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_651
timestamp 1644511149
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_652
timestamp 1644511149
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_653
timestamp 1644511149
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_654
timestamp 1644511149
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_655
timestamp 1644511149
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_656
timestamp 1644511149
transform 1 0 39744 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_657
timestamp 1644511149
transform 1 0 44896 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_658
timestamp 1644511149
transform 1 0 50048 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_659
timestamp 1644511149
transform 1 0 55200 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_660
timestamp 1644511149
transform 1 0 60352 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_661
timestamp 1644511149
transform 1 0 65504 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_662
timestamp 1644511149
transform 1 0 70656 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_663
timestamp 1644511149
transform 1 0 75808 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_664
timestamp 1644511149
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_665
timestamp 1644511149
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_666
timestamp 1644511149
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_667
timestamp 1644511149
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_668
timestamp 1644511149
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_669
timestamp 1644511149
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_670
timestamp 1644511149
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_671
timestamp 1644511149
transform 1 0 42320 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_672
timestamp 1644511149
transform 1 0 47472 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_673
timestamp 1644511149
transform 1 0 52624 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_674
timestamp 1644511149
transform 1 0 57776 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_675
timestamp 1644511149
transform 1 0 62928 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_676
timestamp 1644511149
transform 1 0 68080 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_677
timestamp 1644511149
transform 1 0 73232 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_678
timestamp 1644511149
transform 1 0 78384 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_679
timestamp 1644511149
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_680
timestamp 1644511149
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_681
timestamp 1644511149
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_682
timestamp 1644511149
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_683
timestamp 1644511149
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_684
timestamp 1644511149
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_685
timestamp 1644511149
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_686
timestamp 1644511149
transform 1 0 39744 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_687
timestamp 1644511149
transform 1 0 44896 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_688
timestamp 1644511149
transform 1 0 50048 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_689
timestamp 1644511149
transform 1 0 55200 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_690
timestamp 1644511149
transform 1 0 60352 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_691
timestamp 1644511149
transform 1 0 65504 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_692
timestamp 1644511149
transform 1 0 70656 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_693
timestamp 1644511149
transform 1 0 75808 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_694
timestamp 1644511149
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_695
timestamp 1644511149
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_696
timestamp 1644511149
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_697
timestamp 1644511149
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_698
timestamp 1644511149
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_699
timestamp 1644511149
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_700
timestamp 1644511149
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_701
timestamp 1644511149
transform 1 0 42320 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_702
timestamp 1644511149
transform 1 0 47472 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_703
timestamp 1644511149
transform 1 0 52624 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_704
timestamp 1644511149
transform 1 0 57776 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_705
timestamp 1644511149
transform 1 0 62928 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_706
timestamp 1644511149
transform 1 0 68080 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_707
timestamp 1644511149
transform 1 0 73232 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_708
timestamp 1644511149
transform 1 0 78384 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_709
timestamp 1644511149
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_710
timestamp 1644511149
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_711
timestamp 1644511149
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_712
timestamp 1644511149
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_713
timestamp 1644511149
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_714
timestamp 1644511149
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_715
timestamp 1644511149
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_716
timestamp 1644511149
transform 1 0 39744 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_717
timestamp 1644511149
transform 1 0 44896 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_718
timestamp 1644511149
transform 1 0 50048 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_719
timestamp 1644511149
transform 1 0 55200 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_720
timestamp 1644511149
transform 1 0 60352 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_721
timestamp 1644511149
transform 1 0 65504 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_722
timestamp 1644511149
transform 1 0 70656 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_723
timestamp 1644511149
transform 1 0 75808 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_724
timestamp 1644511149
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_725
timestamp 1644511149
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_726
timestamp 1644511149
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_727
timestamp 1644511149
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_728
timestamp 1644511149
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_729
timestamp 1644511149
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_730
timestamp 1644511149
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_731
timestamp 1644511149
transform 1 0 42320 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_732
timestamp 1644511149
transform 1 0 47472 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_733
timestamp 1644511149
transform 1 0 52624 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_734
timestamp 1644511149
transform 1 0 57776 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_735
timestamp 1644511149
transform 1 0 62928 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_736
timestamp 1644511149
transform 1 0 68080 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_737
timestamp 1644511149
transform 1 0 73232 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_738
timestamp 1644511149
transform 1 0 78384 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_739
timestamp 1644511149
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_740
timestamp 1644511149
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_741
timestamp 1644511149
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_742
timestamp 1644511149
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_743
timestamp 1644511149
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_744
timestamp 1644511149
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_745
timestamp 1644511149
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_746
timestamp 1644511149
transform 1 0 39744 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_747
timestamp 1644511149
transform 1 0 44896 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_748
timestamp 1644511149
transform 1 0 50048 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_749
timestamp 1644511149
transform 1 0 55200 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_750
timestamp 1644511149
transform 1 0 60352 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_751
timestamp 1644511149
transform 1 0 65504 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_752
timestamp 1644511149
transform 1 0 70656 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_753
timestamp 1644511149
transform 1 0 75808 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_754
timestamp 1644511149
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_755
timestamp 1644511149
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_756
timestamp 1644511149
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_757
timestamp 1644511149
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_758
timestamp 1644511149
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_759
timestamp 1644511149
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_760
timestamp 1644511149
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_761
timestamp 1644511149
transform 1 0 42320 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_762
timestamp 1644511149
transform 1 0 47472 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_763
timestamp 1644511149
transform 1 0 52624 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_764
timestamp 1644511149
transform 1 0 57776 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_765
timestamp 1644511149
transform 1 0 62928 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_766
timestamp 1644511149
transform 1 0 68080 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_767
timestamp 1644511149
transform 1 0 73232 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_768
timestamp 1644511149
transform 1 0 78384 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_769
timestamp 1644511149
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_770
timestamp 1644511149
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_771
timestamp 1644511149
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_772
timestamp 1644511149
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_773
timestamp 1644511149
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_774
timestamp 1644511149
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_775
timestamp 1644511149
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_776
timestamp 1644511149
transform 1 0 39744 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_777
timestamp 1644511149
transform 1 0 44896 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_778
timestamp 1644511149
transform 1 0 50048 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_779
timestamp 1644511149
transform 1 0 55200 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_780
timestamp 1644511149
transform 1 0 60352 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_781
timestamp 1644511149
transform 1 0 65504 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_782
timestamp 1644511149
transform 1 0 70656 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_783
timestamp 1644511149
transform 1 0 75808 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_784
timestamp 1644511149
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_785
timestamp 1644511149
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_786
timestamp 1644511149
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_787
timestamp 1644511149
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_788
timestamp 1644511149
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_789
timestamp 1644511149
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_790
timestamp 1644511149
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_791
timestamp 1644511149
transform 1 0 42320 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_792
timestamp 1644511149
transform 1 0 47472 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_793
timestamp 1644511149
transform 1 0 52624 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_794
timestamp 1644511149
transform 1 0 57776 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_795
timestamp 1644511149
transform 1 0 62928 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_796
timestamp 1644511149
transform 1 0 68080 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_797
timestamp 1644511149
transform 1 0 73232 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_798
timestamp 1644511149
transform 1 0 78384 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_799
timestamp 1644511149
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_800
timestamp 1644511149
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_801
timestamp 1644511149
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_802
timestamp 1644511149
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_803
timestamp 1644511149
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_804
timestamp 1644511149
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_805
timestamp 1644511149
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_806
timestamp 1644511149
transform 1 0 39744 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_807
timestamp 1644511149
transform 1 0 44896 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_808
timestamp 1644511149
transform 1 0 50048 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_809
timestamp 1644511149
transform 1 0 55200 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_810
timestamp 1644511149
transform 1 0 60352 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_811
timestamp 1644511149
transform 1 0 65504 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_812
timestamp 1644511149
transform 1 0 70656 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_813
timestamp 1644511149
transform 1 0 75808 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_814
timestamp 1644511149
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_815
timestamp 1644511149
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_816
timestamp 1644511149
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_817
timestamp 1644511149
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_818
timestamp 1644511149
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_819
timestamp 1644511149
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_820
timestamp 1644511149
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_821
timestamp 1644511149
transform 1 0 42320 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_822
timestamp 1644511149
transform 1 0 47472 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_823
timestamp 1644511149
transform 1 0 52624 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_824
timestamp 1644511149
transform 1 0 57776 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_825
timestamp 1644511149
transform 1 0 62928 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_826
timestamp 1644511149
transform 1 0 68080 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_827
timestamp 1644511149
transform 1 0 73232 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_828
timestamp 1644511149
transform 1 0 78384 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_829
timestamp 1644511149
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_830
timestamp 1644511149
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_831
timestamp 1644511149
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_832
timestamp 1644511149
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_833
timestamp 1644511149
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_834
timestamp 1644511149
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_835
timestamp 1644511149
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_836
timestamp 1644511149
transform 1 0 39744 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_837
timestamp 1644511149
transform 1 0 44896 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_838
timestamp 1644511149
transform 1 0 50048 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_839
timestamp 1644511149
transform 1 0 55200 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_840
timestamp 1644511149
transform 1 0 60352 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_841
timestamp 1644511149
transform 1 0 65504 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_842
timestamp 1644511149
transform 1 0 70656 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_843
timestamp 1644511149
transform 1 0 75808 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_844
timestamp 1644511149
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_845
timestamp 1644511149
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_846
timestamp 1644511149
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_847
timestamp 1644511149
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_848
timestamp 1644511149
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_849
timestamp 1644511149
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_850
timestamp 1644511149
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_851
timestamp 1644511149
transform 1 0 42320 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_852
timestamp 1644511149
transform 1 0 47472 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_853
timestamp 1644511149
transform 1 0 52624 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_854
timestamp 1644511149
transform 1 0 57776 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_855
timestamp 1644511149
transform 1 0 62928 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_856
timestamp 1644511149
transform 1 0 68080 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_857
timestamp 1644511149
transform 1 0 73232 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_858
timestamp 1644511149
transform 1 0 78384 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_859
timestamp 1644511149
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_860
timestamp 1644511149
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_861
timestamp 1644511149
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_862
timestamp 1644511149
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_863
timestamp 1644511149
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_864
timestamp 1644511149
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_865
timestamp 1644511149
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_866
timestamp 1644511149
transform 1 0 39744 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_867
timestamp 1644511149
transform 1 0 44896 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_868
timestamp 1644511149
transform 1 0 50048 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_869
timestamp 1644511149
transform 1 0 55200 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_870
timestamp 1644511149
transform 1 0 60352 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_871
timestamp 1644511149
transform 1 0 65504 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_872
timestamp 1644511149
transform 1 0 70656 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_873
timestamp 1644511149
transform 1 0 75808 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_874
timestamp 1644511149
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_875
timestamp 1644511149
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_876
timestamp 1644511149
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_877
timestamp 1644511149
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_878
timestamp 1644511149
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_879
timestamp 1644511149
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_880
timestamp 1644511149
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_881
timestamp 1644511149
transform 1 0 42320 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_882
timestamp 1644511149
transform 1 0 47472 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_883
timestamp 1644511149
transform 1 0 52624 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_884
timestamp 1644511149
transform 1 0 57776 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_885
timestamp 1644511149
transform 1 0 62928 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_886
timestamp 1644511149
transform 1 0 68080 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_887
timestamp 1644511149
transform 1 0 73232 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_888
timestamp 1644511149
transform 1 0 78384 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_889
timestamp 1644511149
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_890
timestamp 1644511149
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_891
timestamp 1644511149
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_892
timestamp 1644511149
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_893
timestamp 1644511149
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_894
timestamp 1644511149
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_895
timestamp 1644511149
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_896
timestamp 1644511149
transform 1 0 39744 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_897
timestamp 1644511149
transform 1 0 44896 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_898
timestamp 1644511149
transform 1 0 50048 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_899
timestamp 1644511149
transform 1 0 55200 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_900
timestamp 1644511149
transform 1 0 60352 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_901
timestamp 1644511149
transform 1 0 65504 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_902
timestamp 1644511149
transform 1 0 70656 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_903
timestamp 1644511149
transform 1 0 75808 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_904
timestamp 1644511149
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_905
timestamp 1644511149
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_906
timestamp 1644511149
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_907
timestamp 1644511149
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_908
timestamp 1644511149
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_909
timestamp 1644511149
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_910
timestamp 1644511149
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_911
timestamp 1644511149
transform 1 0 42320 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_912
timestamp 1644511149
transform 1 0 47472 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_913
timestamp 1644511149
transform 1 0 52624 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_914
timestamp 1644511149
transform 1 0 57776 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_915
timestamp 1644511149
transform 1 0 62928 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_916
timestamp 1644511149
transform 1 0 68080 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_917
timestamp 1644511149
transform 1 0 73232 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_918
timestamp 1644511149
transform 1 0 78384 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_919
timestamp 1644511149
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_920
timestamp 1644511149
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_921
timestamp 1644511149
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_922
timestamp 1644511149
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_923
timestamp 1644511149
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_924
timestamp 1644511149
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_925
timestamp 1644511149
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_926
timestamp 1644511149
transform 1 0 39744 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_927
timestamp 1644511149
transform 1 0 44896 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_928
timestamp 1644511149
transform 1 0 50048 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_929
timestamp 1644511149
transform 1 0 55200 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_930
timestamp 1644511149
transform 1 0 60352 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_931
timestamp 1644511149
transform 1 0 65504 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_932
timestamp 1644511149
transform 1 0 70656 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_933
timestamp 1644511149
transform 1 0 75808 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_934
timestamp 1644511149
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_935
timestamp 1644511149
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_936
timestamp 1644511149
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_937
timestamp 1644511149
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_938
timestamp 1644511149
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_939
timestamp 1644511149
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_940
timestamp 1644511149
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_941
timestamp 1644511149
transform 1 0 42320 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_942
timestamp 1644511149
transform 1 0 47472 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_943
timestamp 1644511149
transform 1 0 52624 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_944
timestamp 1644511149
transform 1 0 57776 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_945
timestamp 1644511149
transform 1 0 62928 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_946
timestamp 1644511149
transform 1 0 68080 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_947
timestamp 1644511149
transform 1 0 73232 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_948
timestamp 1644511149
transform 1 0 78384 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_949
timestamp 1644511149
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_950
timestamp 1644511149
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_951
timestamp 1644511149
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_952
timestamp 1644511149
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_953
timestamp 1644511149
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_954
timestamp 1644511149
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_955
timestamp 1644511149
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_956
timestamp 1644511149
transform 1 0 39744 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_957
timestamp 1644511149
transform 1 0 44896 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_958
timestamp 1644511149
transform 1 0 50048 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_959
timestamp 1644511149
transform 1 0 55200 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_960
timestamp 1644511149
transform 1 0 60352 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_961
timestamp 1644511149
transform 1 0 65504 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_962
timestamp 1644511149
transform 1 0 70656 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_963
timestamp 1644511149
transform 1 0 75808 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_964
timestamp 1644511149
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_965
timestamp 1644511149
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_966
timestamp 1644511149
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_967
timestamp 1644511149
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_968
timestamp 1644511149
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_969
timestamp 1644511149
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_970
timestamp 1644511149
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_971
timestamp 1644511149
transform 1 0 42320 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_972
timestamp 1644511149
transform 1 0 47472 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_973
timestamp 1644511149
transform 1 0 52624 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_974
timestamp 1644511149
transform 1 0 57776 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_975
timestamp 1644511149
transform 1 0 62928 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_976
timestamp 1644511149
transform 1 0 68080 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_977
timestamp 1644511149
transform 1 0 73232 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_978
timestamp 1644511149
transform 1 0 78384 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_979
timestamp 1644511149
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_980
timestamp 1644511149
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_981
timestamp 1644511149
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_982
timestamp 1644511149
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_983
timestamp 1644511149
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_984
timestamp 1644511149
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_985
timestamp 1644511149
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_986
timestamp 1644511149
transform 1 0 39744 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_987
timestamp 1644511149
transform 1 0 44896 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_988
timestamp 1644511149
transform 1 0 50048 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_989
timestamp 1644511149
transform 1 0 55200 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_990
timestamp 1644511149
transform 1 0 60352 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_991
timestamp 1644511149
transform 1 0 65504 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_992
timestamp 1644511149
transform 1 0 70656 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_993
timestamp 1644511149
transform 1 0 75808 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_994
timestamp 1644511149
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_995
timestamp 1644511149
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_996
timestamp 1644511149
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_997
timestamp 1644511149
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_998
timestamp 1644511149
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_999
timestamp 1644511149
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1000
timestamp 1644511149
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1001
timestamp 1644511149
transform 1 0 42320 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1002
timestamp 1644511149
transform 1 0 47472 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1003
timestamp 1644511149
transform 1 0 52624 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1004
timestamp 1644511149
transform 1 0 57776 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1005
timestamp 1644511149
transform 1 0 62928 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1006
timestamp 1644511149
transform 1 0 68080 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1007
timestamp 1644511149
transform 1 0 73232 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1008
timestamp 1644511149
transform 1 0 78384 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1009
timestamp 1644511149
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1010
timestamp 1644511149
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1011
timestamp 1644511149
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1012
timestamp 1644511149
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1013
timestamp 1644511149
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1014
timestamp 1644511149
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1015
timestamp 1644511149
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1016
timestamp 1644511149
transform 1 0 39744 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1017
timestamp 1644511149
transform 1 0 44896 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1018
timestamp 1644511149
transform 1 0 50048 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1019
timestamp 1644511149
transform 1 0 55200 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1020
timestamp 1644511149
transform 1 0 60352 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1021
timestamp 1644511149
transform 1 0 65504 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1022
timestamp 1644511149
transform 1 0 70656 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1023
timestamp 1644511149
transform 1 0 75808 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1024
timestamp 1644511149
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1025
timestamp 1644511149
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1026
timestamp 1644511149
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1027
timestamp 1644511149
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1028
timestamp 1644511149
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1029
timestamp 1644511149
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1030
timestamp 1644511149
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1031
timestamp 1644511149
transform 1 0 42320 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1032
timestamp 1644511149
transform 1 0 47472 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1033
timestamp 1644511149
transform 1 0 52624 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1034
timestamp 1644511149
transform 1 0 57776 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1035
timestamp 1644511149
transform 1 0 62928 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1036
timestamp 1644511149
transform 1 0 68080 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1037
timestamp 1644511149
transform 1 0 73232 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1038
timestamp 1644511149
transform 1 0 78384 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1039
timestamp 1644511149
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1040
timestamp 1644511149
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1041
timestamp 1644511149
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1042
timestamp 1644511149
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1043
timestamp 1644511149
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1044
timestamp 1644511149
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1045
timestamp 1644511149
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1046
timestamp 1644511149
transform 1 0 39744 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1047
timestamp 1644511149
transform 1 0 44896 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1048
timestamp 1644511149
transform 1 0 50048 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1049
timestamp 1644511149
transform 1 0 55200 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1050
timestamp 1644511149
transform 1 0 60352 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1051
timestamp 1644511149
transform 1 0 65504 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1052
timestamp 1644511149
transform 1 0 70656 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1053
timestamp 1644511149
transform 1 0 75808 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1054
timestamp 1644511149
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1055
timestamp 1644511149
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1056
timestamp 1644511149
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1057
timestamp 1644511149
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1058
timestamp 1644511149
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1059
timestamp 1644511149
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1060
timestamp 1644511149
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1061
timestamp 1644511149
transform 1 0 42320 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1062
timestamp 1644511149
transform 1 0 47472 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1063
timestamp 1644511149
transform 1 0 52624 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1064
timestamp 1644511149
transform 1 0 57776 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1065
timestamp 1644511149
transform 1 0 62928 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1066
timestamp 1644511149
transform 1 0 68080 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1067
timestamp 1644511149
transform 1 0 73232 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1068
timestamp 1644511149
transform 1 0 78384 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1069
timestamp 1644511149
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1070
timestamp 1644511149
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1071
timestamp 1644511149
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1072
timestamp 1644511149
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1073
timestamp 1644511149
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1074
timestamp 1644511149
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1075
timestamp 1644511149
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1076
timestamp 1644511149
transform 1 0 39744 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1077
timestamp 1644511149
transform 1 0 44896 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1078
timestamp 1644511149
transform 1 0 50048 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1079
timestamp 1644511149
transform 1 0 55200 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1080
timestamp 1644511149
transform 1 0 60352 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1081
timestamp 1644511149
transform 1 0 65504 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1082
timestamp 1644511149
transform 1 0 70656 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1083
timestamp 1644511149
transform 1 0 75808 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1084
timestamp 1644511149
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1085
timestamp 1644511149
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1086
timestamp 1644511149
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1087
timestamp 1644511149
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1088
timestamp 1644511149
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1089
timestamp 1644511149
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1090
timestamp 1644511149
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1091
timestamp 1644511149
transform 1 0 42320 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1092
timestamp 1644511149
transform 1 0 47472 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1093
timestamp 1644511149
transform 1 0 52624 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1094
timestamp 1644511149
transform 1 0 57776 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1095
timestamp 1644511149
transform 1 0 62928 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1096
timestamp 1644511149
transform 1 0 68080 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1097
timestamp 1644511149
transform 1 0 73232 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1098
timestamp 1644511149
transform 1 0 78384 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1099
timestamp 1644511149
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1100
timestamp 1644511149
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1101
timestamp 1644511149
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1102
timestamp 1644511149
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1103
timestamp 1644511149
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1104
timestamp 1644511149
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1105
timestamp 1644511149
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1106
timestamp 1644511149
transform 1 0 39744 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1107
timestamp 1644511149
transform 1 0 44896 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1108
timestamp 1644511149
transform 1 0 50048 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1109
timestamp 1644511149
transform 1 0 55200 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1110
timestamp 1644511149
transform 1 0 60352 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1111
timestamp 1644511149
transform 1 0 65504 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1112
timestamp 1644511149
transform 1 0 70656 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1113
timestamp 1644511149
transform 1 0 75808 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1114
timestamp 1644511149
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1115
timestamp 1644511149
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1116
timestamp 1644511149
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1117
timestamp 1644511149
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1118
timestamp 1644511149
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1119
timestamp 1644511149
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1120
timestamp 1644511149
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1121
timestamp 1644511149
transform 1 0 42320 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1122
timestamp 1644511149
transform 1 0 47472 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1123
timestamp 1644511149
transform 1 0 52624 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1124
timestamp 1644511149
transform 1 0 57776 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1125
timestamp 1644511149
transform 1 0 62928 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1126
timestamp 1644511149
transform 1 0 68080 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1127
timestamp 1644511149
transform 1 0 73232 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1128
timestamp 1644511149
transform 1 0 78384 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1129
timestamp 1644511149
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1130
timestamp 1644511149
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1131
timestamp 1644511149
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1132
timestamp 1644511149
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1133
timestamp 1644511149
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1134
timestamp 1644511149
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1135
timestamp 1644511149
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1136
timestamp 1644511149
transform 1 0 39744 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1137
timestamp 1644511149
transform 1 0 44896 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1138
timestamp 1644511149
transform 1 0 50048 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1139
timestamp 1644511149
transform 1 0 55200 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1140
timestamp 1644511149
transform 1 0 60352 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1141
timestamp 1644511149
transform 1 0 65504 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1142
timestamp 1644511149
transform 1 0 70656 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1143
timestamp 1644511149
transform 1 0 75808 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1144
timestamp 1644511149
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1145
timestamp 1644511149
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1146
timestamp 1644511149
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1147
timestamp 1644511149
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1148
timestamp 1644511149
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1149
timestamp 1644511149
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1150
timestamp 1644511149
transform 1 0 37168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1151
timestamp 1644511149
transform 1 0 42320 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1152
timestamp 1644511149
transform 1 0 47472 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1153
timestamp 1644511149
transform 1 0 52624 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1154
timestamp 1644511149
transform 1 0 57776 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1155
timestamp 1644511149
transform 1 0 62928 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1156
timestamp 1644511149
transform 1 0 68080 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1157
timestamp 1644511149
transform 1 0 73232 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1158
timestamp 1644511149
transform 1 0 78384 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1159
timestamp 1644511149
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1160
timestamp 1644511149
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1161
timestamp 1644511149
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1162
timestamp 1644511149
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1163
timestamp 1644511149
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1164
timestamp 1644511149
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1165
timestamp 1644511149
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1166
timestamp 1644511149
transform 1 0 39744 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1167
timestamp 1644511149
transform 1 0 44896 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1168
timestamp 1644511149
transform 1 0 50048 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1169
timestamp 1644511149
transform 1 0 55200 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1170
timestamp 1644511149
transform 1 0 60352 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1171
timestamp 1644511149
transform 1 0 65504 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1172
timestamp 1644511149
transform 1 0 70656 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1173
timestamp 1644511149
transform 1 0 75808 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1174
timestamp 1644511149
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1175
timestamp 1644511149
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1176
timestamp 1644511149
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1177
timestamp 1644511149
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1178
timestamp 1644511149
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1179
timestamp 1644511149
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1180
timestamp 1644511149
transform 1 0 37168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1181
timestamp 1644511149
transform 1 0 42320 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1182
timestamp 1644511149
transform 1 0 47472 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1183
timestamp 1644511149
transform 1 0 52624 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1184
timestamp 1644511149
transform 1 0 57776 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1185
timestamp 1644511149
transform 1 0 62928 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1186
timestamp 1644511149
transform 1 0 68080 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1187
timestamp 1644511149
transform 1 0 73232 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1188
timestamp 1644511149
transform 1 0 78384 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1189
timestamp 1644511149
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1190
timestamp 1644511149
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1191
timestamp 1644511149
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1192
timestamp 1644511149
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1193
timestamp 1644511149
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1194
timestamp 1644511149
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1195
timestamp 1644511149
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1196
timestamp 1644511149
transform 1 0 39744 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1197
timestamp 1644511149
transform 1 0 44896 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1198
timestamp 1644511149
transform 1 0 50048 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1199
timestamp 1644511149
transform 1 0 55200 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1200
timestamp 1644511149
transform 1 0 60352 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1201
timestamp 1644511149
transform 1 0 65504 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1202
timestamp 1644511149
transform 1 0 70656 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1203
timestamp 1644511149
transform 1 0 75808 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1204
timestamp 1644511149
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1205
timestamp 1644511149
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1206
timestamp 1644511149
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1207
timestamp 1644511149
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1208
timestamp 1644511149
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1209
timestamp 1644511149
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1210
timestamp 1644511149
transform 1 0 37168 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1211
timestamp 1644511149
transform 1 0 42320 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1212
timestamp 1644511149
transform 1 0 47472 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1213
timestamp 1644511149
transform 1 0 52624 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1214
timestamp 1644511149
transform 1 0 57776 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1215
timestamp 1644511149
transform 1 0 62928 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1216
timestamp 1644511149
transform 1 0 68080 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1217
timestamp 1644511149
transform 1 0 73232 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1218
timestamp 1644511149
transform 1 0 78384 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1219
timestamp 1644511149
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1220
timestamp 1644511149
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1221
timestamp 1644511149
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1222
timestamp 1644511149
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1223
timestamp 1644511149
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1224
timestamp 1644511149
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1225
timestamp 1644511149
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1226
timestamp 1644511149
transform 1 0 39744 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1227
timestamp 1644511149
transform 1 0 44896 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1228
timestamp 1644511149
transform 1 0 50048 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1229
timestamp 1644511149
transform 1 0 55200 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1230
timestamp 1644511149
transform 1 0 60352 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1231
timestamp 1644511149
transform 1 0 65504 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1232
timestamp 1644511149
transform 1 0 70656 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1233
timestamp 1644511149
transform 1 0 75808 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1234
timestamp 1644511149
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1235
timestamp 1644511149
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1236
timestamp 1644511149
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1237
timestamp 1644511149
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1238
timestamp 1644511149
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1239
timestamp 1644511149
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1240
timestamp 1644511149
transform 1 0 37168 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1241
timestamp 1644511149
transform 1 0 42320 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1242
timestamp 1644511149
transform 1 0 47472 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1243
timestamp 1644511149
transform 1 0 52624 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1244
timestamp 1644511149
transform 1 0 57776 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1245
timestamp 1644511149
transform 1 0 62928 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1246
timestamp 1644511149
transform 1 0 68080 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1247
timestamp 1644511149
transform 1 0 73232 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1248
timestamp 1644511149
transform 1 0 78384 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1249
timestamp 1644511149
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1250
timestamp 1644511149
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1251
timestamp 1644511149
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1252
timestamp 1644511149
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1253
timestamp 1644511149
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1254
timestamp 1644511149
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1255
timestamp 1644511149
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1256
timestamp 1644511149
transform 1 0 39744 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1257
timestamp 1644511149
transform 1 0 44896 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1258
timestamp 1644511149
transform 1 0 50048 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1259
timestamp 1644511149
transform 1 0 55200 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1260
timestamp 1644511149
transform 1 0 60352 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1261
timestamp 1644511149
transform 1 0 65504 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1262
timestamp 1644511149
transform 1 0 70656 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1263
timestamp 1644511149
transform 1 0 75808 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1264
timestamp 1644511149
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1265
timestamp 1644511149
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1266
timestamp 1644511149
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1267
timestamp 1644511149
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1268
timestamp 1644511149
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1269
timestamp 1644511149
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1270
timestamp 1644511149
transform 1 0 37168 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1271
timestamp 1644511149
transform 1 0 42320 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1272
timestamp 1644511149
transform 1 0 47472 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1273
timestamp 1644511149
transform 1 0 52624 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1274
timestamp 1644511149
transform 1 0 57776 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1275
timestamp 1644511149
transform 1 0 62928 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1276
timestamp 1644511149
transform 1 0 68080 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1277
timestamp 1644511149
transform 1 0 73232 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1278
timestamp 1644511149
transform 1 0 78384 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1279
timestamp 1644511149
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1280
timestamp 1644511149
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1281
timestamp 1644511149
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1282
timestamp 1644511149
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1283
timestamp 1644511149
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1284
timestamp 1644511149
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1285
timestamp 1644511149
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1286
timestamp 1644511149
transform 1 0 39744 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1287
timestamp 1644511149
transform 1 0 44896 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1288
timestamp 1644511149
transform 1 0 50048 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1289
timestamp 1644511149
transform 1 0 55200 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1290
timestamp 1644511149
transform 1 0 60352 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1291
timestamp 1644511149
transform 1 0 65504 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1292
timestamp 1644511149
transform 1 0 70656 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1293
timestamp 1644511149
transform 1 0 75808 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1294
timestamp 1644511149
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1295
timestamp 1644511149
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1296
timestamp 1644511149
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1297
timestamp 1644511149
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1298
timestamp 1644511149
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1299
timestamp 1644511149
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1300
timestamp 1644511149
transform 1 0 37168 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1301
timestamp 1644511149
transform 1 0 42320 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1302
timestamp 1644511149
transform 1 0 47472 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1303
timestamp 1644511149
transform 1 0 52624 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1304
timestamp 1644511149
transform 1 0 57776 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1305
timestamp 1644511149
transform 1 0 62928 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1306
timestamp 1644511149
transform 1 0 68080 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1307
timestamp 1644511149
transform 1 0 73232 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1308
timestamp 1644511149
transform 1 0 78384 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1309
timestamp 1644511149
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1310
timestamp 1644511149
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1311
timestamp 1644511149
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1312
timestamp 1644511149
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1313
timestamp 1644511149
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1314
timestamp 1644511149
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1315
timestamp 1644511149
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1316
timestamp 1644511149
transform 1 0 39744 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1317
timestamp 1644511149
transform 1 0 44896 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1318
timestamp 1644511149
transform 1 0 50048 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1319
timestamp 1644511149
transform 1 0 55200 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1320
timestamp 1644511149
transform 1 0 60352 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1321
timestamp 1644511149
transform 1 0 65504 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1322
timestamp 1644511149
transform 1 0 70656 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1323
timestamp 1644511149
transform 1 0 75808 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1324
timestamp 1644511149
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1325
timestamp 1644511149
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1326
timestamp 1644511149
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1327
timestamp 1644511149
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1328
timestamp 1644511149
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1329
timestamp 1644511149
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1330
timestamp 1644511149
transform 1 0 37168 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1331
timestamp 1644511149
transform 1 0 42320 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1332
timestamp 1644511149
transform 1 0 47472 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1333
timestamp 1644511149
transform 1 0 52624 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1334
timestamp 1644511149
transform 1 0 57776 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1335
timestamp 1644511149
transform 1 0 62928 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1336
timestamp 1644511149
transform 1 0 68080 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1337
timestamp 1644511149
transform 1 0 73232 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1338
timestamp 1644511149
transform 1 0 78384 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1339
timestamp 1644511149
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1340
timestamp 1644511149
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1341
timestamp 1644511149
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1342
timestamp 1644511149
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1343
timestamp 1644511149
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1344
timestamp 1644511149
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1345
timestamp 1644511149
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1346
timestamp 1644511149
transform 1 0 39744 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1347
timestamp 1644511149
transform 1 0 44896 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1348
timestamp 1644511149
transform 1 0 50048 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1349
timestamp 1644511149
transform 1 0 55200 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1350
timestamp 1644511149
transform 1 0 60352 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1351
timestamp 1644511149
transform 1 0 65504 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1352
timestamp 1644511149
transform 1 0 70656 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1353
timestamp 1644511149
transform 1 0 75808 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1354
timestamp 1644511149
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1355
timestamp 1644511149
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1356
timestamp 1644511149
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1357
timestamp 1644511149
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1358
timestamp 1644511149
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1359
timestamp 1644511149
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1360
timestamp 1644511149
transform 1 0 37168 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1361
timestamp 1644511149
transform 1 0 42320 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1362
timestamp 1644511149
transform 1 0 47472 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1363
timestamp 1644511149
transform 1 0 52624 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1364
timestamp 1644511149
transform 1 0 57776 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1365
timestamp 1644511149
transform 1 0 62928 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1366
timestamp 1644511149
transform 1 0 68080 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1367
timestamp 1644511149
transform 1 0 73232 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1368
timestamp 1644511149
transform 1 0 78384 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1369
timestamp 1644511149
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1370
timestamp 1644511149
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1371
timestamp 1644511149
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1372
timestamp 1644511149
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1373
timestamp 1644511149
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1374
timestamp 1644511149
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1375
timestamp 1644511149
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1376
timestamp 1644511149
transform 1 0 39744 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1377
timestamp 1644511149
transform 1 0 44896 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1378
timestamp 1644511149
transform 1 0 50048 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1379
timestamp 1644511149
transform 1 0 55200 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1380
timestamp 1644511149
transform 1 0 60352 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1381
timestamp 1644511149
transform 1 0 65504 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1382
timestamp 1644511149
transform 1 0 70656 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1383
timestamp 1644511149
transform 1 0 75808 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1384
timestamp 1644511149
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1385
timestamp 1644511149
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1386
timestamp 1644511149
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1387
timestamp 1644511149
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1388
timestamp 1644511149
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1389
timestamp 1644511149
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1390
timestamp 1644511149
transform 1 0 37168 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1391
timestamp 1644511149
transform 1 0 42320 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1392
timestamp 1644511149
transform 1 0 47472 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1393
timestamp 1644511149
transform 1 0 52624 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1394
timestamp 1644511149
transform 1 0 57776 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1395
timestamp 1644511149
transform 1 0 62928 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1396
timestamp 1644511149
transform 1 0 68080 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1397
timestamp 1644511149
transform 1 0 73232 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1398
timestamp 1644511149
transform 1 0 78384 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1399
timestamp 1644511149
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1400
timestamp 1644511149
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1401
timestamp 1644511149
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1402
timestamp 1644511149
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1403
timestamp 1644511149
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1404
timestamp 1644511149
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1405
timestamp 1644511149
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1406
timestamp 1644511149
transform 1 0 39744 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1407
timestamp 1644511149
transform 1 0 44896 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1408
timestamp 1644511149
transform 1 0 50048 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1409
timestamp 1644511149
transform 1 0 55200 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1410
timestamp 1644511149
transform 1 0 60352 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1411
timestamp 1644511149
transform 1 0 65504 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1412
timestamp 1644511149
transform 1 0 70656 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1413
timestamp 1644511149
transform 1 0 75808 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1414
timestamp 1644511149
transform 1 0 6256 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1415
timestamp 1644511149
transform 1 0 11408 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1416
timestamp 1644511149
transform 1 0 16560 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1417
timestamp 1644511149
transform 1 0 21712 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1418
timestamp 1644511149
transform 1 0 26864 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1419
timestamp 1644511149
transform 1 0 32016 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1420
timestamp 1644511149
transform 1 0 37168 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1421
timestamp 1644511149
transform 1 0 42320 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1422
timestamp 1644511149
transform 1 0 47472 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1423
timestamp 1644511149
transform 1 0 52624 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1424
timestamp 1644511149
transform 1 0 57776 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1425
timestamp 1644511149
transform 1 0 62928 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1426
timestamp 1644511149
transform 1 0 68080 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1427
timestamp 1644511149
transform 1 0 73232 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1428
timestamp 1644511149
transform 1 0 78384 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1429
timestamp 1644511149
transform 1 0 3680 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1430
timestamp 1644511149
transform 1 0 8832 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1431
timestamp 1644511149
transform 1 0 13984 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1432
timestamp 1644511149
transform 1 0 19136 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1433
timestamp 1644511149
transform 1 0 24288 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1434
timestamp 1644511149
transform 1 0 29440 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1435
timestamp 1644511149
transform 1 0 34592 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1436
timestamp 1644511149
transform 1 0 39744 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1437
timestamp 1644511149
transform 1 0 44896 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1438
timestamp 1644511149
transform 1 0 50048 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1439
timestamp 1644511149
transform 1 0 55200 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1440
timestamp 1644511149
transform 1 0 60352 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1441
timestamp 1644511149
transform 1 0 65504 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1442
timestamp 1644511149
transform 1 0 70656 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1443
timestamp 1644511149
transform 1 0 75808 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1444
timestamp 1644511149
transform 1 0 6256 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1445
timestamp 1644511149
transform 1 0 11408 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1446
timestamp 1644511149
transform 1 0 16560 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1447
timestamp 1644511149
transform 1 0 21712 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1448
timestamp 1644511149
transform 1 0 26864 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1449
timestamp 1644511149
transform 1 0 32016 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1450
timestamp 1644511149
transform 1 0 37168 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1451
timestamp 1644511149
transform 1 0 42320 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1452
timestamp 1644511149
transform 1 0 47472 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1453
timestamp 1644511149
transform 1 0 52624 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1454
timestamp 1644511149
transform 1 0 57776 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1455
timestamp 1644511149
transform 1 0 62928 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1456
timestamp 1644511149
transform 1 0 68080 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1457
timestamp 1644511149
transform 1 0 73232 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1458
timestamp 1644511149
transform 1 0 78384 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1459
timestamp 1644511149
transform 1 0 3680 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1460
timestamp 1644511149
transform 1 0 8832 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1461
timestamp 1644511149
transform 1 0 13984 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1462
timestamp 1644511149
transform 1 0 19136 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1463
timestamp 1644511149
transform 1 0 24288 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1464
timestamp 1644511149
transform 1 0 29440 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1465
timestamp 1644511149
transform 1 0 34592 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1466
timestamp 1644511149
transform 1 0 39744 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1467
timestamp 1644511149
transform 1 0 44896 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1468
timestamp 1644511149
transform 1 0 50048 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1469
timestamp 1644511149
transform 1 0 55200 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1470
timestamp 1644511149
transform 1 0 60352 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1471
timestamp 1644511149
transform 1 0 65504 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1472
timestamp 1644511149
transform 1 0 70656 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1473
timestamp 1644511149
transform 1 0 75808 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1474
timestamp 1644511149
transform 1 0 6256 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1475
timestamp 1644511149
transform 1 0 11408 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1476
timestamp 1644511149
transform 1 0 16560 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1477
timestamp 1644511149
transform 1 0 21712 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1478
timestamp 1644511149
transform 1 0 26864 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1479
timestamp 1644511149
transform 1 0 32016 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1480
timestamp 1644511149
transform 1 0 37168 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1481
timestamp 1644511149
transform 1 0 42320 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1482
timestamp 1644511149
transform 1 0 47472 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1483
timestamp 1644511149
transform 1 0 52624 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1484
timestamp 1644511149
transform 1 0 57776 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1485
timestamp 1644511149
transform 1 0 62928 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1486
timestamp 1644511149
transform 1 0 68080 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1487
timestamp 1644511149
transform 1 0 73232 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1488
timestamp 1644511149
transform 1 0 78384 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1489
timestamp 1644511149
transform 1 0 3680 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1490
timestamp 1644511149
transform 1 0 8832 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1491
timestamp 1644511149
transform 1 0 13984 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1492
timestamp 1644511149
transform 1 0 19136 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1493
timestamp 1644511149
transform 1 0 24288 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1494
timestamp 1644511149
transform 1 0 29440 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1495
timestamp 1644511149
transform 1 0 34592 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1496
timestamp 1644511149
transform 1 0 39744 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1497
timestamp 1644511149
transform 1 0 44896 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1498
timestamp 1644511149
transform 1 0 50048 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1499
timestamp 1644511149
transform 1 0 55200 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1500
timestamp 1644511149
transform 1 0 60352 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1501
timestamp 1644511149
transform 1 0 65504 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1502
timestamp 1644511149
transform 1 0 70656 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1503
timestamp 1644511149
transform 1 0 75808 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1504
timestamp 1644511149
transform 1 0 6256 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1505
timestamp 1644511149
transform 1 0 11408 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1506
timestamp 1644511149
transform 1 0 16560 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1507
timestamp 1644511149
transform 1 0 21712 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1508
timestamp 1644511149
transform 1 0 26864 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1509
timestamp 1644511149
transform 1 0 32016 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1510
timestamp 1644511149
transform 1 0 37168 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1511
timestamp 1644511149
transform 1 0 42320 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1512
timestamp 1644511149
transform 1 0 47472 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1513
timestamp 1644511149
transform 1 0 52624 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1514
timestamp 1644511149
transform 1 0 57776 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1515
timestamp 1644511149
transform 1 0 62928 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1516
timestamp 1644511149
transform 1 0 68080 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1517
timestamp 1644511149
transform 1 0 73232 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1518
timestamp 1644511149
transform 1 0 78384 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1519
timestamp 1644511149
transform 1 0 3680 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1520
timestamp 1644511149
transform 1 0 8832 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1521
timestamp 1644511149
transform 1 0 13984 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1522
timestamp 1644511149
transform 1 0 19136 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1523
timestamp 1644511149
transform 1 0 24288 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1524
timestamp 1644511149
transform 1 0 29440 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1525
timestamp 1644511149
transform 1 0 34592 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1526
timestamp 1644511149
transform 1 0 39744 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1527
timestamp 1644511149
transform 1 0 44896 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1528
timestamp 1644511149
transform 1 0 50048 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1529
timestamp 1644511149
transform 1 0 55200 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1530
timestamp 1644511149
transform 1 0 60352 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1531
timestamp 1644511149
transform 1 0 65504 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1532
timestamp 1644511149
transform 1 0 70656 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1533
timestamp 1644511149
transform 1 0 75808 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1534
timestamp 1644511149
transform 1 0 6256 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1535
timestamp 1644511149
transform 1 0 11408 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1536
timestamp 1644511149
transform 1 0 16560 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1537
timestamp 1644511149
transform 1 0 21712 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1538
timestamp 1644511149
transform 1 0 26864 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1539
timestamp 1644511149
transform 1 0 32016 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1540
timestamp 1644511149
transform 1 0 37168 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1541
timestamp 1644511149
transform 1 0 42320 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1542
timestamp 1644511149
transform 1 0 47472 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1543
timestamp 1644511149
transform 1 0 52624 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1544
timestamp 1644511149
transform 1 0 57776 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1545
timestamp 1644511149
transform 1 0 62928 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1546
timestamp 1644511149
transform 1 0 68080 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1547
timestamp 1644511149
transform 1 0 73232 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1548
timestamp 1644511149
transform 1 0 78384 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1549
timestamp 1644511149
transform 1 0 3680 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1550
timestamp 1644511149
transform 1 0 8832 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1551
timestamp 1644511149
transform 1 0 13984 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1552
timestamp 1644511149
transform 1 0 19136 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1553
timestamp 1644511149
transform 1 0 24288 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1554
timestamp 1644511149
transform 1 0 29440 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1555
timestamp 1644511149
transform 1 0 34592 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1556
timestamp 1644511149
transform 1 0 39744 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1557
timestamp 1644511149
transform 1 0 44896 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1558
timestamp 1644511149
transform 1 0 50048 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1559
timestamp 1644511149
transform 1 0 55200 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1560
timestamp 1644511149
transform 1 0 60352 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1561
timestamp 1644511149
transform 1 0 65504 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1562
timestamp 1644511149
transform 1 0 70656 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1563
timestamp 1644511149
transform 1 0 75808 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1564
timestamp 1644511149
transform 1 0 6256 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1565
timestamp 1644511149
transform 1 0 11408 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1566
timestamp 1644511149
transform 1 0 16560 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1567
timestamp 1644511149
transform 1 0 21712 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1568
timestamp 1644511149
transform 1 0 26864 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1569
timestamp 1644511149
transform 1 0 32016 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1570
timestamp 1644511149
transform 1 0 37168 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1571
timestamp 1644511149
transform 1 0 42320 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1572
timestamp 1644511149
transform 1 0 47472 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1573
timestamp 1644511149
transform 1 0 52624 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1574
timestamp 1644511149
transform 1 0 57776 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1575
timestamp 1644511149
transform 1 0 62928 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1576
timestamp 1644511149
transform 1 0 68080 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1577
timestamp 1644511149
transform 1 0 73232 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1578
timestamp 1644511149
transform 1 0 78384 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1579
timestamp 1644511149
transform 1 0 3680 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1580
timestamp 1644511149
transform 1 0 8832 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1581
timestamp 1644511149
transform 1 0 13984 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1582
timestamp 1644511149
transform 1 0 19136 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1583
timestamp 1644511149
transform 1 0 24288 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1584
timestamp 1644511149
transform 1 0 29440 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1585
timestamp 1644511149
transform 1 0 34592 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1586
timestamp 1644511149
transform 1 0 39744 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1587
timestamp 1644511149
transform 1 0 44896 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1588
timestamp 1644511149
transform 1 0 50048 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1589
timestamp 1644511149
transform 1 0 55200 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1590
timestamp 1644511149
transform 1 0 60352 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1591
timestamp 1644511149
transform 1 0 65504 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1592
timestamp 1644511149
transform 1 0 70656 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1593
timestamp 1644511149
transform 1 0 75808 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1594
timestamp 1644511149
transform 1 0 6256 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1595
timestamp 1644511149
transform 1 0 11408 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1596
timestamp 1644511149
transform 1 0 16560 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1597
timestamp 1644511149
transform 1 0 21712 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1598
timestamp 1644511149
transform 1 0 26864 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1599
timestamp 1644511149
transform 1 0 32016 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1600
timestamp 1644511149
transform 1 0 37168 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1601
timestamp 1644511149
transform 1 0 42320 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1602
timestamp 1644511149
transform 1 0 47472 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1603
timestamp 1644511149
transform 1 0 52624 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1604
timestamp 1644511149
transform 1 0 57776 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1605
timestamp 1644511149
transform 1 0 62928 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1606
timestamp 1644511149
transform 1 0 68080 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1607
timestamp 1644511149
transform 1 0 73232 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1608
timestamp 1644511149
transform 1 0 78384 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1609
timestamp 1644511149
transform 1 0 3680 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1610
timestamp 1644511149
transform 1 0 8832 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1611
timestamp 1644511149
transform 1 0 13984 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1612
timestamp 1644511149
transform 1 0 19136 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1613
timestamp 1644511149
transform 1 0 24288 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1614
timestamp 1644511149
transform 1 0 29440 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1615
timestamp 1644511149
transform 1 0 34592 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1616
timestamp 1644511149
transform 1 0 39744 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1617
timestamp 1644511149
transform 1 0 44896 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1618
timestamp 1644511149
transform 1 0 50048 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1619
timestamp 1644511149
transform 1 0 55200 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1620
timestamp 1644511149
transform 1 0 60352 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1621
timestamp 1644511149
transform 1 0 65504 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1622
timestamp 1644511149
transform 1 0 70656 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1623
timestamp 1644511149
transform 1 0 75808 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1624
timestamp 1644511149
transform 1 0 6256 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1625
timestamp 1644511149
transform 1 0 11408 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1626
timestamp 1644511149
transform 1 0 16560 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1627
timestamp 1644511149
transform 1 0 21712 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1628
timestamp 1644511149
transform 1 0 26864 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1629
timestamp 1644511149
transform 1 0 32016 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1630
timestamp 1644511149
transform 1 0 37168 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1631
timestamp 1644511149
transform 1 0 42320 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1632
timestamp 1644511149
transform 1 0 47472 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1633
timestamp 1644511149
transform 1 0 52624 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1634
timestamp 1644511149
transform 1 0 57776 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1635
timestamp 1644511149
transform 1 0 62928 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1636
timestamp 1644511149
transform 1 0 68080 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1637
timestamp 1644511149
transform 1 0 73232 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1638
timestamp 1644511149
transform 1 0 78384 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1639
timestamp 1644511149
transform 1 0 3680 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1640
timestamp 1644511149
transform 1 0 8832 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1641
timestamp 1644511149
transform 1 0 13984 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1642
timestamp 1644511149
transform 1 0 19136 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1643
timestamp 1644511149
transform 1 0 24288 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1644
timestamp 1644511149
transform 1 0 29440 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1645
timestamp 1644511149
transform 1 0 34592 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1646
timestamp 1644511149
transform 1 0 39744 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1647
timestamp 1644511149
transform 1 0 44896 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1648
timestamp 1644511149
transform 1 0 50048 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1649
timestamp 1644511149
transform 1 0 55200 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1650
timestamp 1644511149
transform 1 0 60352 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1651
timestamp 1644511149
transform 1 0 65504 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1652
timestamp 1644511149
transform 1 0 70656 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1653
timestamp 1644511149
transform 1 0 75808 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1654
timestamp 1644511149
transform 1 0 6256 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1655
timestamp 1644511149
transform 1 0 11408 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1656
timestamp 1644511149
transform 1 0 16560 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1657
timestamp 1644511149
transform 1 0 21712 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1658
timestamp 1644511149
transform 1 0 26864 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1659
timestamp 1644511149
transform 1 0 32016 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1660
timestamp 1644511149
transform 1 0 37168 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1661
timestamp 1644511149
transform 1 0 42320 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1662
timestamp 1644511149
transform 1 0 47472 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1663
timestamp 1644511149
transform 1 0 52624 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1664
timestamp 1644511149
transform 1 0 57776 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1665
timestamp 1644511149
transform 1 0 62928 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1666
timestamp 1644511149
transform 1 0 68080 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1667
timestamp 1644511149
transform 1 0 73232 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1668
timestamp 1644511149
transform 1 0 78384 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1669
timestamp 1644511149
transform 1 0 3680 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1670
timestamp 1644511149
transform 1 0 8832 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1671
timestamp 1644511149
transform 1 0 13984 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1672
timestamp 1644511149
transform 1 0 19136 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1673
timestamp 1644511149
transform 1 0 24288 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1674
timestamp 1644511149
transform 1 0 29440 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1675
timestamp 1644511149
transform 1 0 34592 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1676
timestamp 1644511149
transform 1 0 39744 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1677
timestamp 1644511149
transform 1 0 44896 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1678
timestamp 1644511149
transform 1 0 50048 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1679
timestamp 1644511149
transform 1 0 55200 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1680
timestamp 1644511149
transform 1 0 60352 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1681
timestamp 1644511149
transform 1 0 65504 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1682
timestamp 1644511149
transform 1 0 70656 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1683
timestamp 1644511149
transform 1 0 75808 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1684
timestamp 1644511149
transform 1 0 6256 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1685
timestamp 1644511149
transform 1 0 11408 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1686
timestamp 1644511149
transform 1 0 16560 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1687
timestamp 1644511149
transform 1 0 21712 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1688
timestamp 1644511149
transform 1 0 26864 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1689
timestamp 1644511149
transform 1 0 32016 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1690
timestamp 1644511149
transform 1 0 37168 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1691
timestamp 1644511149
transform 1 0 42320 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1692
timestamp 1644511149
transform 1 0 47472 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1693
timestamp 1644511149
transform 1 0 52624 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1694
timestamp 1644511149
transform 1 0 57776 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1695
timestamp 1644511149
transform 1 0 62928 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1696
timestamp 1644511149
transform 1 0 68080 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1697
timestamp 1644511149
transform 1 0 73232 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1698
timestamp 1644511149
transform 1 0 78384 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1699
timestamp 1644511149
transform 1 0 3680 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1700
timestamp 1644511149
transform 1 0 8832 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1701
timestamp 1644511149
transform 1 0 13984 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1702
timestamp 1644511149
transform 1 0 19136 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1703
timestamp 1644511149
transform 1 0 24288 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1704
timestamp 1644511149
transform 1 0 29440 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1705
timestamp 1644511149
transform 1 0 34592 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1706
timestamp 1644511149
transform 1 0 39744 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1707
timestamp 1644511149
transform 1 0 44896 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1708
timestamp 1644511149
transform 1 0 50048 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1709
timestamp 1644511149
transform 1 0 55200 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1710
timestamp 1644511149
transform 1 0 60352 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1711
timestamp 1644511149
transform 1 0 65504 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1712
timestamp 1644511149
transform 1 0 70656 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1713
timestamp 1644511149
transform 1 0 75808 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1714
timestamp 1644511149
transform 1 0 6256 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1715
timestamp 1644511149
transform 1 0 11408 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1716
timestamp 1644511149
transform 1 0 16560 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1717
timestamp 1644511149
transform 1 0 21712 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1718
timestamp 1644511149
transform 1 0 26864 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1719
timestamp 1644511149
transform 1 0 32016 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1720
timestamp 1644511149
transform 1 0 37168 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1721
timestamp 1644511149
transform 1 0 42320 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1722
timestamp 1644511149
transform 1 0 47472 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1723
timestamp 1644511149
transform 1 0 52624 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1724
timestamp 1644511149
transform 1 0 57776 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1725
timestamp 1644511149
transform 1 0 62928 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1726
timestamp 1644511149
transform 1 0 68080 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1727
timestamp 1644511149
transform 1 0 73232 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1728
timestamp 1644511149
transform 1 0 78384 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1729
timestamp 1644511149
transform 1 0 3680 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1730
timestamp 1644511149
transform 1 0 8832 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1731
timestamp 1644511149
transform 1 0 13984 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1732
timestamp 1644511149
transform 1 0 19136 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1733
timestamp 1644511149
transform 1 0 24288 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1734
timestamp 1644511149
transform 1 0 29440 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1735
timestamp 1644511149
transform 1 0 34592 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1736
timestamp 1644511149
transform 1 0 39744 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1737
timestamp 1644511149
transform 1 0 44896 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1738
timestamp 1644511149
transform 1 0 50048 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1739
timestamp 1644511149
transform 1 0 55200 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1740
timestamp 1644511149
transform 1 0 60352 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1741
timestamp 1644511149
transform 1 0 65504 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1742
timestamp 1644511149
transform 1 0 70656 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1743
timestamp 1644511149
transform 1 0 75808 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1744
timestamp 1644511149
transform 1 0 6256 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1745
timestamp 1644511149
transform 1 0 11408 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1746
timestamp 1644511149
transform 1 0 16560 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1747
timestamp 1644511149
transform 1 0 21712 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1748
timestamp 1644511149
transform 1 0 26864 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1749
timestamp 1644511149
transform 1 0 32016 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1750
timestamp 1644511149
transform 1 0 37168 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1751
timestamp 1644511149
transform 1 0 42320 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1752
timestamp 1644511149
transform 1 0 47472 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1753
timestamp 1644511149
transform 1 0 52624 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1754
timestamp 1644511149
transform 1 0 57776 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1755
timestamp 1644511149
transform 1 0 62928 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1756
timestamp 1644511149
transform 1 0 68080 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1757
timestamp 1644511149
transform 1 0 73232 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1758
timestamp 1644511149
transform 1 0 78384 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1759
timestamp 1644511149
transform 1 0 3680 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1760
timestamp 1644511149
transform 1 0 8832 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1761
timestamp 1644511149
transform 1 0 13984 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1762
timestamp 1644511149
transform 1 0 19136 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1763
timestamp 1644511149
transform 1 0 24288 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1764
timestamp 1644511149
transform 1 0 29440 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1765
timestamp 1644511149
transform 1 0 34592 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1766
timestamp 1644511149
transform 1 0 39744 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1767
timestamp 1644511149
transform 1 0 44896 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1768
timestamp 1644511149
transform 1 0 50048 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1769
timestamp 1644511149
transform 1 0 55200 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1770
timestamp 1644511149
transform 1 0 60352 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1771
timestamp 1644511149
transform 1 0 65504 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1772
timestamp 1644511149
transform 1 0 70656 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1773
timestamp 1644511149
transform 1 0 75808 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1774
timestamp 1644511149
transform 1 0 6256 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1775
timestamp 1644511149
transform 1 0 11408 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1776
timestamp 1644511149
transform 1 0 16560 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1777
timestamp 1644511149
transform 1 0 21712 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1778
timestamp 1644511149
transform 1 0 26864 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1779
timestamp 1644511149
transform 1 0 32016 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1780
timestamp 1644511149
transform 1 0 37168 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1781
timestamp 1644511149
transform 1 0 42320 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1782
timestamp 1644511149
transform 1 0 47472 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1783
timestamp 1644511149
transform 1 0 52624 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1784
timestamp 1644511149
transform 1 0 57776 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1785
timestamp 1644511149
transform 1 0 62928 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1786
timestamp 1644511149
transform 1 0 68080 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1787
timestamp 1644511149
transform 1 0 73232 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1788
timestamp 1644511149
transform 1 0 78384 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1789
timestamp 1644511149
transform 1 0 3680 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1790
timestamp 1644511149
transform 1 0 8832 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1791
timestamp 1644511149
transform 1 0 13984 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1792
timestamp 1644511149
transform 1 0 19136 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1793
timestamp 1644511149
transform 1 0 24288 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1794
timestamp 1644511149
transform 1 0 29440 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1795
timestamp 1644511149
transform 1 0 34592 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1796
timestamp 1644511149
transform 1 0 39744 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1797
timestamp 1644511149
transform 1 0 44896 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1798
timestamp 1644511149
transform 1 0 50048 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1799
timestamp 1644511149
transform 1 0 55200 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1800
timestamp 1644511149
transform 1 0 60352 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1801
timestamp 1644511149
transform 1 0 65504 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1802
timestamp 1644511149
transform 1 0 70656 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1803
timestamp 1644511149
transform 1 0 75808 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1804
timestamp 1644511149
transform 1 0 6256 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1805
timestamp 1644511149
transform 1 0 11408 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1806
timestamp 1644511149
transform 1 0 16560 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1807
timestamp 1644511149
transform 1 0 21712 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1808
timestamp 1644511149
transform 1 0 26864 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1809
timestamp 1644511149
transform 1 0 32016 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1810
timestamp 1644511149
transform 1 0 37168 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1811
timestamp 1644511149
transform 1 0 42320 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1812
timestamp 1644511149
transform 1 0 47472 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1813
timestamp 1644511149
transform 1 0 52624 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1814
timestamp 1644511149
transform 1 0 57776 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1815
timestamp 1644511149
transform 1 0 62928 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1816
timestamp 1644511149
transform 1 0 68080 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1817
timestamp 1644511149
transform 1 0 73232 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1818
timestamp 1644511149
transform 1 0 78384 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1819
timestamp 1644511149
transform 1 0 3680 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1820
timestamp 1644511149
transform 1 0 8832 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1821
timestamp 1644511149
transform 1 0 13984 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1822
timestamp 1644511149
transform 1 0 19136 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1823
timestamp 1644511149
transform 1 0 24288 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1824
timestamp 1644511149
transform 1 0 29440 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1825
timestamp 1644511149
transform 1 0 34592 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1826
timestamp 1644511149
transform 1 0 39744 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1827
timestamp 1644511149
transform 1 0 44896 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1828
timestamp 1644511149
transform 1 0 50048 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1829
timestamp 1644511149
transform 1 0 55200 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1830
timestamp 1644511149
transform 1 0 60352 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1831
timestamp 1644511149
transform 1 0 65504 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1832
timestamp 1644511149
transform 1 0 70656 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1833
timestamp 1644511149
transform 1 0 75808 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1834
timestamp 1644511149
transform 1 0 6256 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1835
timestamp 1644511149
transform 1 0 11408 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1836
timestamp 1644511149
transform 1 0 16560 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1837
timestamp 1644511149
transform 1 0 21712 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1838
timestamp 1644511149
transform 1 0 26864 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1839
timestamp 1644511149
transform 1 0 32016 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1840
timestamp 1644511149
transform 1 0 37168 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1841
timestamp 1644511149
transform 1 0 42320 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1842
timestamp 1644511149
transform 1 0 47472 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1843
timestamp 1644511149
transform 1 0 52624 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1844
timestamp 1644511149
transform 1 0 57776 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1845
timestamp 1644511149
transform 1 0 62928 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1846
timestamp 1644511149
transform 1 0 68080 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1847
timestamp 1644511149
transform 1 0 73232 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1848
timestamp 1644511149
transform 1 0 78384 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1849
timestamp 1644511149
transform 1 0 3680 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1850
timestamp 1644511149
transform 1 0 8832 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1851
timestamp 1644511149
transform 1 0 13984 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1852
timestamp 1644511149
transform 1 0 19136 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1853
timestamp 1644511149
transform 1 0 24288 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1854
timestamp 1644511149
transform 1 0 29440 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1855
timestamp 1644511149
transform 1 0 34592 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1856
timestamp 1644511149
transform 1 0 39744 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1857
timestamp 1644511149
transform 1 0 44896 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1858
timestamp 1644511149
transform 1 0 50048 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1859
timestamp 1644511149
transform 1 0 55200 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1860
timestamp 1644511149
transform 1 0 60352 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1861
timestamp 1644511149
transform 1 0 65504 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1862
timestamp 1644511149
transform 1 0 70656 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1863
timestamp 1644511149
transform 1 0 75808 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1864
timestamp 1644511149
transform 1 0 6256 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1865
timestamp 1644511149
transform 1 0 11408 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1866
timestamp 1644511149
transform 1 0 16560 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1867
timestamp 1644511149
transform 1 0 21712 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1868
timestamp 1644511149
transform 1 0 26864 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1869
timestamp 1644511149
transform 1 0 32016 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1870
timestamp 1644511149
transform 1 0 37168 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1871
timestamp 1644511149
transform 1 0 42320 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1872
timestamp 1644511149
transform 1 0 47472 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1873
timestamp 1644511149
transform 1 0 52624 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1874
timestamp 1644511149
transform 1 0 57776 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1875
timestamp 1644511149
transform 1 0 62928 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1876
timestamp 1644511149
transform 1 0 68080 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1877
timestamp 1644511149
transform 1 0 73232 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1878
timestamp 1644511149
transform 1 0 78384 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1879
timestamp 1644511149
transform 1 0 3680 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1880
timestamp 1644511149
transform 1 0 8832 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1881
timestamp 1644511149
transform 1 0 13984 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1882
timestamp 1644511149
transform 1 0 19136 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1883
timestamp 1644511149
transform 1 0 24288 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1884
timestamp 1644511149
transform 1 0 29440 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1885
timestamp 1644511149
transform 1 0 34592 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1886
timestamp 1644511149
transform 1 0 39744 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1887
timestamp 1644511149
transform 1 0 44896 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1888
timestamp 1644511149
transform 1 0 50048 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1889
timestamp 1644511149
transform 1 0 55200 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1890
timestamp 1644511149
transform 1 0 60352 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1891
timestamp 1644511149
transform 1 0 65504 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1892
timestamp 1644511149
transform 1 0 70656 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1893
timestamp 1644511149
transform 1 0 75808 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1894
timestamp 1644511149
transform 1 0 6256 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1895
timestamp 1644511149
transform 1 0 11408 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1896
timestamp 1644511149
transform 1 0 16560 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1897
timestamp 1644511149
transform 1 0 21712 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1898
timestamp 1644511149
transform 1 0 26864 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1899
timestamp 1644511149
transform 1 0 32016 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1900
timestamp 1644511149
transform 1 0 37168 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1901
timestamp 1644511149
transform 1 0 42320 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1902
timestamp 1644511149
transform 1 0 47472 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1903
timestamp 1644511149
transform 1 0 52624 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1904
timestamp 1644511149
transform 1 0 57776 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1905
timestamp 1644511149
transform 1 0 62928 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1906
timestamp 1644511149
transform 1 0 68080 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1907
timestamp 1644511149
transform 1 0 73232 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1908
timestamp 1644511149
transform 1 0 78384 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1909
timestamp 1644511149
transform 1 0 3680 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1910
timestamp 1644511149
transform 1 0 8832 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1911
timestamp 1644511149
transform 1 0 13984 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1912
timestamp 1644511149
transform 1 0 19136 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1913
timestamp 1644511149
transform 1 0 24288 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1914
timestamp 1644511149
transform 1 0 29440 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1915
timestamp 1644511149
transform 1 0 34592 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1916
timestamp 1644511149
transform 1 0 39744 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1917
timestamp 1644511149
transform 1 0 44896 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1918
timestamp 1644511149
transform 1 0 50048 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1919
timestamp 1644511149
transform 1 0 55200 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1920
timestamp 1644511149
transform 1 0 60352 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1921
timestamp 1644511149
transform 1 0 65504 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1922
timestamp 1644511149
transform 1 0 70656 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1923
timestamp 1644511149
transform 1 0 75808 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1924
timestamp 1644511149
transform 1 0 6256 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1925
timestamp 1644511149
transform 1 0 11408 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1926
timestamp 1644511149
transform 1 0 16560 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1927
timestamp 1644511149
transform 1 0 21712 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1928
timestamp 1644511149
transform 1 0 26864 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1929
timestamp 1644511149
transform 1 0 32016 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1930
timestamp 1644511149
transform 1 0 37168 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1931
timestamp 1644511149
transform 1 0 42320 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1932
timestamp 1644511149
transform 1 0 47472 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1933
timestamp 1644511149
transform 1 0 52624 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1934
timestamp 1644511149
transform 1 0 57776 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1935
timestamp 1644511149
transform 1 0 62928 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1936
timestamp 1644511149
transform 1 0 68080 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1937
timestamp 1644511149
transform 1 0 73232 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1938
timestamp 1644511149
transform 1 0 78384 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1939
timestamp 1644511149
transform 1 0 3680 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1940
timestamp 1644511149
transform 1 0 8832 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1941
timestamp 1644511149
transform 1 0 13984 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1942
timestamp 1644511149
transform 1 0 19136 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1943
timestamp 1644511149
transform 1 0 24288 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1944
timestamp 1644511149
transform 1 0 29440 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1945
timestamp 1644511149
transform 1 0 34592 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1946
timestamp 1644511149
transform 1 0 39744 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1947
timestamp 1644511149
transform 1 0 44896 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1948
timestamp 1644511149
transform 1 0 50048 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1949
timestamp 1644511149
transform 1 0 55200 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1950
timestamp 1644511149
transform 1 0 60352 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1951
timestamp 1644511149
transform 1 0 65504 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1952
timestamp 1644511149
transform 1 0 70656 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1953
timestamp 1644511149
transform 1 0 75808 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1954
timestamp 1644511149
transform 1 0 6256 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1955
timestamp 1644511149
transform 1 0 11408 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1956
timestamp 1644511149
transform 1 0 16560 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1957
timestamp 1644511149
transform 1 0 21712 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1958
timestamp 1644511149
transform 1 0 26864 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1959
timestamp 1644511149
transform 1 0 32016 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1960
timestamp 1644511149
transform 1 0 37168 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1961
timestamp 1644511149
transform 1 0 42320 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1962
timestamp 1644511149
transform 1 0 47472 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1963
timestamp 1644511149
transform 1 0 52624 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1964
timestamp 1644511149
transform 1 0 57776 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1965
timestamp 1644511149
transform 1 0 62928 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1966
timestamp 1644511149
transform 1 0 68080 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1967
timestamp 1644511149
transform 1 0 73232 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1968
timestamp 1644511149
transform 1 0 78384 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1969
timestamp 1644511149
transform 1 0 3680 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1970
timestamp 1644511149
transform 1 0 8832 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1971
timestamp 1644511149
transform 1 0 13984 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1972
timestamp 1644511149
transform 1 0 19136 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1973
timestamp 1644511149
transform 1 0 24288 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1974
timestamp 1644511149
transform 1 0 29440 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1975
timestamp 1644511149
transform 1 0 34592 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1976
timestamp 1644511149
transform 1 0 39744 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1977
timestamp 1644511149
transform 1 0 44896 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1978
timestamp 1644511149
transform 1 0 50048 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1979
timestamp 1644511149
transform 1 0 55200 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1980
timestamp 1644511149
transform 1 0 60352 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1981
timestamp 1644511149
transform 1 0 65504 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1982
timestamp 1644511149
transform 1 0 70656 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1983
timestamp 1644511149
transform 1 0 75808 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1984
timestamp 1644511149
transform 1 0 6256 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1985
timestamp 1644511149
transform 1 0 11408 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1986
timestamp 1644511149
transform 1 0 16560 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1987
timestamp 1644511149
transform 1 0 21712 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1988
timestamp 1644511149
transform 1 0 26864 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1989
timestamp 1644511149
transform 1 0 32016 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1990
timestamp 1644511149
transform 1 0 37168 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1991
timestamp 1644511149
transform 1 0 42320 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1992
timestamp 1644511149
transform 1 0 47472 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1993
timestamp 1644511149
transform 1 0 52624 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1994
timestamp 1644511149
transform 1 0 57776 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1995
timestamp 1644511149
transform 1 0 62928 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1996
timestamp 1644511149
transform 1 0 68080 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1997
timestamp 1644511149
transform 1 0 73232 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1998
timestamp 1644511149
transform 1 0 78384 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1999
timestamp 1644511149
transform 1 0 3680 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2000
timestamp 1644511149
transform 1 0 8832 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2001
timestamp 1644511149
transform 1 0 13984 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2002
timestamp 1644511149
transform 1 0 19136 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2003
timestamp 1644511149
transform 1 0 24288 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2004
timestamp 1644511149
transform 1 0 29440 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2005
timestamp 1644511149
transform 1 0 34592 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2006
timestamp 1644511149
transform 1 0 39744 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2007
timestamp 1644511149
transform 1 0 44896 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2008
timestamp 1644511149
transform 1 0 50048 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2009
timestamp 1644511149
transform 1 0 55200 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2010
timestamp 1644511149
transform 1 0 60352 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2011
timestamp 1644511149
transform 1 0 65504 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2012
timestamp 1644511149
transform 1 0 70656 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2013
timestamp 1644511149
transform 1 0 75808 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2014
timestamp 1644511149
transform 1 0 6256 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2015
timestamp 1644511149
transform 1 0 11408 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2016
timestamp 1644511149
transform 1 0 16560 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2017
timestamp 1644511149
transform 1 0 21712 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2018
timestamp 1644511149
transform 1 0 26864 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2019
timestamp 1644511149
transform 1 0 32016 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2020
timestamp 1644511149
transform 1 0 37168 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2021
timestamp 1644511149
transform 1 0 42320 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2022
timestamp 1644511149
transform 1 0 47472 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2023
timestamp 1644511149
transform 1 0 52624 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2024
timestamp 1644511149
transform 1 0 57776 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2025
timestamp 1644511149
transform 1 0 62928 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2026
timestamp 1644511149
transform 1 0 68080 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2027
timestamp 1644511149
transform 1 0 73232 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2028
timestamp 1644511149
transform 1 0 78384 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2029
timestamp 1644511149
transform 1 0 3680 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2030
timestamp 1644511149
transform 1 0 8832 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2031
timestamp 1644511149
transform 1 0 13984 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2032
timestamp 1644511149
transform 1 0 19136 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2033
timestamp 1644511149
transform 1 0 24288 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2034
timestamp 1644511149
transform 1 0 29440 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2035
timestamp 1644511149
transform 1 0 34592 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2036
timestamp 1644511149
transform 1 0 39744 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2037
timestamp 1644511149
transform 1 0 44896 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2038
timestamp 1644511149
transform 1 0 50048 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2039
timestamp 1644511149
transform 1 0 55200 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2040
timestamp 1644511149
transform 1 0 60352 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2041
timestamp 1644511149
transform 1 0 65504 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2042
timestamp 1644511149
transform 1 0 70656 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2043
timestamp 1644511149
transform 1 0 75808 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2044
timestamp 1644511149
transform 1 0 6256 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2045
timestamp 1644511149
transform 1 0 11408 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2046
timestamp 1644511149
transform 1 0 16560 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2047
timestamp 1644511149
transform 1 0 21712 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2048
timestamp 1644511149
transform 1 0 26864 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2049
timestamp 1644511149
transform 1 0 32016 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2050
timestamp 1644511149
transform 1 0 37168 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2051
timestamp 1644511149
transform 1 0 42320 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2052
timestamp 1644511149
transform 1 0 47472 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2053
timestamp 1644511149
transform 1 0 52624 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2054
timestamp 1644511149
transform 1 0 57776 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2055
timestamp 1644511149
transform 1 0 62928 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2056
timestamp 1644511149
transform 1 0 68080 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2057
timestamp 1644511149
transform 1 0 73232 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2058
timestamp 1644511149
transform 1 0 78384 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2059
timestamp 1644511149
transform 1 0 3680 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2060
timestamp 1644511149
transform 1 0 8832 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2061
timestamp 1644511149
transform 1 0 13984 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2062
timestamp 1644511149
transform 1 0 19136 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2063
timestamp 1644511149
transform 1 0 24288 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2064
timestamp 1644511149
transform 1 0 29440 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2065
timestamp 1644511149
transform 1 0 34592 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2066
timestamp 1644511149
transform 1 0 39744 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2067
timestamp 1644511149
transform 1 0 44896 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2068
timestamp 1644511149
transform 1 0 50048 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2069
timestamp 1644511149
transform 1 0 55200 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2070
timestamp 1644511149
transform 1 0 60352 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2071
timestamp 1644511149
transform 1 0 65504 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2072
timestamp 1644511149
transform 1 0 70656 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2073
timestamp 1644511149
transform 1 0 75808 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2074
timestamp 1644511149
transform 1 0 6256 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2075
timestamp 1644511149
transform 1 0 11408 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2076
timestamp 1644511149
transform 1 0 16560 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2077
timestamp 1644511149
transform 1 0 21712 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2078
timestamp 1644511149
transform 1 0 26864 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2079
timestamp 1644511149
transform 1 0 32016 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2080
timestamp 1644511149
transform 1 0 37168 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2081
timestamp 1644511149
transform 1 0 42320 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2082
timestamp 1644511149
transform 1 0 47472 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2083
timestamp 1644511149
transform 1 0 52624 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2084
timestamp 1644511149
transform 1 0 57776 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2085
timestamp 1644511149
transform 1 0 62928 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2086
timestamp 1644511149
transform 1 0 68080 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2087
timestamp 1644511149
transform 1 0 73232 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2088
timestamp 1644511149
transform 1 0 78384 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2089
timestamp 1644511149
transform 1 0 3680 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2090
timestamp 1644511149
transform 1 0 8832 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2091
timestamp 1644511149
transform 1 0 13984 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2092
timestamp 1644511149
transform 1 0 19136 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2093
timestamp 1644511149
transform 1 0 24288 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2094
timestamp 1644511149
transform 1 0 29440 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2095
timestamp 1644511149
transform 1 0 34592 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2096
timestamp 1644511149
transform 1 0 39744 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2097
timestamp 1644511149
transform 1 0 44896 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2098
timestamp 1644511149
transform 1 0 50048 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2099
timestamp 1644511149
transform 1 0 55200 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2100
timestamp 1644511149
transform 1 0 60352 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2101
timestamp 1644511149
transform 1 0 65504 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2102
timestamp 1644511149
transform 1 0 70656 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2103
timestamp 1644511149
transform 1 0 75808 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2104
timestamp 1644511149
transform 1 0 6256 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2105
timestamp 1644511149
transform 1 0 11408 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2106
timestamp 1644511149
transform 1 0 16560 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2107
timestamp 1644511149
transform 1 0 21712 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2108
timestamp 1644511149
transform 1 0 26864 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2109
timestamp 1644511149
transform 1 0 32016 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2110
timestamp 1644511149
transform 1 0 37168 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2111
timestamp 1644511149
transform 1 0 42320 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2112
timestamp 1644511149
transform 1 0 47472 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2113
timestamp 1644511149
transform 1 0 52624 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2114
timestamp 1644511149
transform 1 0 57776 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2115
timestamp 1644511149
transform 1 0 62928 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2116
timestamp 1644511149
transform 1 0 68080 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2117
timestamp 1644511149
transform 1 0 73232 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2118
timestamp 1644511149
transform 1 0 78384 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2119
timestamp 1644511149
transform 1 0 3680 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2120
timestamp 1644511149
transform 1 0 8832 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2121
timestamp 1644511149
transform 1 0 13984 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2122
timestamp 1644511149
transform 1 0 19136 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2123
timestamp 1644511149
transform 1 0 24288 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2124
timestamp 1644511149
transform 1 0 29440 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2125
timestamp 1644511149
transform 1 0 34592 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2126
timestamp 1644511149
transform 1 0 39744 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2127
timestamp 1644511149
transform 1 0 44896 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2128
timestamp 1644511149
transform 1 0 50048 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2129
timestamp 1644511149
transform 1 0 55200 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2130
timestamp 1644511149
transform 1 0 60352 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2131
timestamp 1644511149
transform 1 0 65504 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2132
timestamp 1644511149
transform 1 0 70656 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2133
timestamp 1644511149
transform 1 0 75808 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2134
timestamp 1644511149
transform 1 0 6256 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2135
timestamp 1644511149
transform 1 0 11408 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2136
timestamp 1644511149
transform 1 0 16560 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2137
timestamp 1644511149
transform 1 0 21712 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2138
timestamp 1644511149
transform 1 0 26864 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2139
timestamp 1644511149
transform 1 0 32016 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2140
timestamp 1644511149
transform 1 0 37168 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2141
timestamp 1644511149
transform 1 0 42320 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2142
timestamp 1644511149
transform 1 0 47472 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2143
timestamp 1644511149
transform 1 0 52624 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2144
timestamp 1644511149
transform 1 0 57776 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2145
timestamp 1644511149
transform 1 0 62928 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2146
timestamp 1644511149
transform 1 0 68080 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2147
timestamp 1644511149
transform 1 0 73232 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2148
timestamp 1644511149
transform 1 0 78384 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2149
timestamp 1644511149
transform 1 0 3680 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2150
timestamp 1644511149
transform 1 0 8832 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2151
timestamp 1644511149
transform 1 0 13984 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2152
timestamp 1644511149
transform 1 0 19136 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2153
timestamp 1644511149
transform 1 0 24288 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2154
timestamp 1644511149
transform 1 0 29440 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2155
timestamp 1644511149
transform 1 0 34592 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2156
timestamp 1644511149
transform 1 0 39744 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2157
timestamp 1644511149
transform 1 0 44896 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2158
timestamp 1644511149
transform 1 0 50048 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2159
timestamp 1644511149
transform 1 0 55200 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2160
timestamp 1644511149
transform 1 0 60352 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2161
timestamp 1644511149
transform 1 0 65504 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2162
timestamp 1644511149
transform 1 0 70656 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2163
timestamp 1644511149
transform 1 0 75808 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2164
timestamp 1644511149
transform 1 0 6256 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2165
timestamp 1644511149
transform 1 0 11408 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2166
timestamp 1644511149
transform 1 0 16560 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2167
timestamp 1644511149
transform 1 0 21712 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2168
timestamp 1644511149
transform 1 0 26864 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2169
timestamp 1644511149
transform 1 0 32016 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2170
timestamp 1644511149
transform 1 0 37168 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2171
timestamp 1644511149
transform 1 0 42320 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2172
timestamp 1644511149
transform 1 0 47472 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2173
timestamp 1644511149
transform 1 0 52624 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2174
timestamp 1644511149
transform 1 0 57776 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2175
timestamp 1644511149
transform 1 0 62928 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2176
timestamp 1644511149
transform 1 0 68080 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2177
timestamp 1644511149
transform 1 0 73232 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2178
timestamp 1644511149
transform 1 0 78384 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2179
timestamp 1644511149
transform 1 0 3680 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2180
timestamp 1644511149
transform 1 0 8832 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2181
timestamp 1644511149
transform 1 0 13984 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2182
timestamp 1644511149
transform 1 0 19136 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2183
timestamp 1644511149
transform 1 0 24288 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2184
timestamp 1644511149
transform 1 0 29440 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2185
timestamp 1644511149
transform 1 0 34592 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2186
timestamp 1644511149
transform 1 0 39744 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2187
timestamp 1644511149
transform 1 0 44896 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2188
timestamp 1644511149
transform 1 0 50048 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2189
timestamp 1644511149
transform 1 0 55200 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2190
timestamp 1644511149
transform 1 0 60352 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2191
timestamp 1644511149
transform 1 0 65504 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2192
timestamp 1644511149
transform 1 0 70656 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2193
timestamp 1644511149
transform 1 0 75808 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2194
timestamp 1644511149
transform 1 0 6256 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2195
timestamp 1644511149
transform 1 0 11408 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2196
timestamp 1644511149
transform 1 0 16560 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2197
timestamp 1644511149
transform 1 0 21712 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2198
timestamp 1644511149
transform 1 0 26864 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2199
timestamp 1644511149
transform 1 0 32016 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2200
timestamp 1644511149
transform 1 0 37168 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2201
timestamp 1644511149
transform 1 0 42320 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2202
timestamp 1644511149
transform 1 0 47472 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2203
timestamp 1644511149
transform 1 0 52624 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2204
timestamp 1644511149
transform 1 0 57776 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2205
timestamp 1644511149
transform 1 0 62928 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2206
timestamp 1644511149
transform 1 0 68080 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2207
timestamp 1644511149
transform 1 0 73232 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2208
timestamp 1644511149
transform 1 0 78384 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2209
timestamp 1644511149
transform 1 0 3680 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2210
timestamp 1644511149
transform 1 0 8832 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2211
timestamp 1644511149
transform 1 0 13984 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2212
timestamp 1644511149
transform 1 0 19136 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2213
timestamp 1644511149
transform 1 0 24288 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2214
timestamp 1644511149
transform 1 0 29440 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2215
timestamp 1644511149
transform 1 0 34592 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2216
timestamp 1644511149
transform 1 0 39744 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2217
timestamp 1644511149
transform 1 0 44896 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2218
timestamp 1644511149
transform 1 0 50048 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2219
timestamp 1644511149
transform 1 0 55200 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2220
timestamp 1644511149
transform 1 0 60352 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2221
timestamp 1644511149
transform 1 0 65504 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2222
timestamp 1644511149
transform 1 0 70656 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2223
timestamp 1644511149
transform 1 0 75808 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2224
timestamp 1644511149
transform 1 0 6256 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2225
timestamp 1644511149
transform 1 0 11408 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2226
timestamp 1644511149
transform 1 0 16560 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2227
timestamp 1644511149
transform 1 0 21712 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2228
timestamp 1644511149
transform 1 0 26864 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2229
timestamp 1644511149
transform 1 0 32016 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2230
timestamp 1644511149
transform 1 0 37168 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2231
timestamp 1644511149
transform 1 0 42320 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2232
timestamp 1644511149
transform 1 0 47472 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2233
timestamp 1644511149
transform 1 0 52624 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2234
timestamp 1644511149
transform 1 0 57776 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2235
timestamp 1644511149
transform 1 0 62928 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2236
timestamp 1644511149
transform 1 0 68080 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2237
timestamp 1644511149
transform 1 0 73232 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2238
timestamp 1644511149
transform 1 0 78384 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2239
timestamp 1644511149
transform 1 0 3680 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2240
timestamp 1644511149
transform 1 0 8832 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2241
timestamp 1644511149
transform 1 0 13984 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2242
timestamp 1644511149
transform 1 0 19136 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2243
timestamp 1644511149
transform 1 0 24288 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2244
timestamp 1644511149
transform 1 0 29440 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2245
timestamp 1644511149
transform 1 0 34592 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2246
timestamp 1644511149
transform 1 0 39744 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2247
timestamp 1644511149
transform 1 0 44896 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2248
timestamp 1644511149
transform 1 0 50048 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2249
timestamp 1644511149
transform 1 0 55200 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2250
timestamp 1644511149
transform 1 0 60352 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2251
timestamp 1644511149
transform 1 0 65504 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2252
timestamp 1644511149
transform 1 0 70656 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2253
timestamp 1644511149
transform 1 0 75808 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2254
timestamp 1644511149
transform 1 0 6256 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2255
timestamp 1644511149
transform 1 0 11408 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2256
timestamp 1644511149
transform 1 0 16560 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2257
timestamp 1644511149
transform 1 0 21712 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2258
timestamp 1644511149
transform 1 0 26864 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2259
timestamp 1644511149
transform 1 0 32016 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2260
timestamp 1644511149
transform 1 0 37168 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2261
timestamp 1644511149
transform 1 0 42320 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2262
timestamp 1644511149
transform 1 0 47472 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2263
timestamp 1644511149
transform 1 0 52624 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2264
timestamp 1644511149
transform 1 0 57776 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2265
timestamp 1644511149
transform 1 0 62928 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2266
timestamp 1644511149
transform 1 0 68080 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2267
timestamp 1644511149
transform 1 0 73232 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2268
timestamp 1644511149
transform 1 0 78384 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2269
timestamp 1644511149
transform 1 0 3680 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2270
timestamp 1644511149
transform 1 0 8832 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2271
timestamp 1644511149
transform 1 0 13984 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2272
timestamp 1644511149
transform 1 0 19136 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2273
timestamp 1644511149
transform 1 0 24288 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2274
timestamp 1644511149
transform 1 0 29440 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2275
timestamp 1644511149
transform 1 0 34592 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2276
timestamp 1644511149
transform 1 0 39744 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2277
timestamp 1644511149
transform 1 0 44896 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2278
timestamp 1644511149
transform 1 0 50048 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2279
timestamp 1644511149
transform 1 0 55200 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2280
timestamp 1644511149
transform 1 0 60352 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2281
timestamp 1644511149
transform 1 0 65504 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2282
timestamp 1644511149
transform 1 0 70656 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2283
timestamp 1644511149
transform 1 0 75808 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2284
timestamp 1644511149
transform 1 0 6256 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2285
timestamp 1644511149
transform 1 0 11408 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2286
timestamp 1644511149
transform 1 0 16560 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2287
timestamp 1644511149
transform 1 0 21712 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2288
timestamp 1644511149
transform 1 0 26864 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2289
timestamp 1644511149
transform 1 0 32016 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2290
timestamp 1644511149
transform 1 0 37168 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2291
timestamp 1644511149
transform 1 0 42320 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2292
timestamp 1644511149
transform 1 0 47472 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2293
timestamp 1644511149
transform 1 0 52624 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2294
timestamp 1644511149
transform 1 0 57776 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2295
timestamp 1644511149
transform 1 0 62928 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2296
timestamp 1644511149
transform 1 0 68080 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2297
timestamp 1644511149
transform 1 0 73232 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2298
timestamp 1644511149
transform 1 0 78384 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2299
timestamp 1644511149
transform 1 0 3680 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2300
timestamp 1644511149
transform 1 0 8832 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2301
timestamp 1644511149
transform 1 0 13984 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2302
timestamp 1644511149
transform 1 0 19136 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2303
timestamp 1644511149
transform 1 0 24288 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2304
timestamp 1644511149
transform 1 0 29440 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2305
timestamp 1644511149
transform 1 0 34592 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2306
timestamp 1644511149
transform 1 0 39744 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2307
timestamp 1644511149
transform 1 0 44896 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2308
timestamp 1644511149
transform 1 0 50048 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2309
timestamp 1644511149
transform 1 0 55200 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2310
timestamp 1644511149
transform 1 0 60352 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2311
timestamp 1644511149
transform 1 0 65504 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2312
timestamp 1644511149
transform 1 0 70656 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2313
timestamp 1644511149
transform 1 0 75808 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2314
timestamp 1644511149
transform 1 0 6256 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2315
timestamp 1644511149
transform 1 0 11408 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2316
timestamp 1644511149
transform 1 0 16560 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2317
timestamp 1644511149
transform 1 0 21712 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2318
timestamp 1644511149
transform 1 0 26864 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2319
timestamp 1644511149
transform 1 0 32016 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2320
timestamp 1644511149
transform 1 0 37168 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2321
timestamp 1644511149
transform 1 0 42320 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2322
timestamp 1644511149
transform 1 0 47472 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2323
timestamp 1644511149
transform 1 0 52624 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2324
timestamp 1644511149
transform 1 0 57776 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2325
timestamp 1644511149
transform 1 0 62928 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2326
timestamp 1644511149
transform 1 0 68080 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2327
timestamp 1644511149
transform 1 0 73232 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2328
timestamp 1644511149
transform 1 0 78384 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2329
timestamp 1644511149
transform 1 0 3680 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2330
timestamp 1644511149
transform 1 0 8832 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2331
timestamp 1644511149
transform 1 0 13984 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2332
timestamp 1644511149
transform 1 0 19136 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2333
timestamp 1644511149
transform 1 0 24288 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2334
timestamp 1644511149
transform 1 0 29440 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2335
timestamp 1644511149
transform 1 0 34592 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2336
timestamp 1644511149
transform 1 0 39744 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2337
timestamp 1644511149
transform 1 0 44896 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2338
timestamp 1644511149
transform 1 0 50048 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2339
timestamp 1644511149
transform 1 0 55200 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2340
timestamp 1644511149
transform 1 0 60352 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2341
timestamp 1644511149
transform 1 0 65504 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2342
timestamp 1644511149
transform 1 0 70656 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2343
timestamp 1644511149
transform 1 0 75808 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2344
timestamp 1644511149
transform 1 0 6256 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2345
timestamp 1644511149
transform 1 0 11408 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2346
timestamp 1644511149
transform 1 0 16560 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2347
timestamp 1644511149
transform 1 0 21712 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2348
timestamp 1644511149
transform 1 0 26864 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2349
timestamp 1644511149
transform 1 0 32016 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2350
timestamp 1644511149
transform 1 0 37168 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2351
timestamp 1644511149
transform 1 0 42320 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2352
timestamp 1644511149
transform 1 0 47472 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2353
timestamp 1644511149
transform 1 0 52624 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2354
timestamp 1644511149
transform 1 0 57776 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2355
timestamp 1644511149
transform 1 0 62928 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2356
timestamp 1644511149
transform 1 0 68080 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2357
timestamp 1644511149
transform 1 0 73232 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2358
timestamp 1644511149
transform 1 0 78384 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2359
timestamp 1644511149
transform 1 0 3680 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2360
timestamp 1644511149
transform 1 0 8832 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2361
timestamp 1644511149
transform 1 0 13984 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2362
timestamp 1644511149
transform 1 0 19136 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2363
timestamp 1644511149
transform 1 0 24288 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2364
timestamp 1644511149
transform 1 0 29440 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2365
timestamp 1644511149
transform 1 0 34592 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2366
timestamp 1644511149
transform 1 0 39744 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2367
timestamp 1644511149
transform 1 0 44896 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2368
timestamp 1644511149
transform 1 0 50048 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2369
timestamp 1644511149
transform 1 0 55200 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2370
timestamp 1644511149
transform 1 0 60352 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2371
timestamp 1644511149
transform 1 0 65504 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2372
timestamp 1644511149
transform 1 0 70656 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2373
timestamp 1644511149
transform 1 0 75808 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2374
timestamp 1644511149
transform 1 0 6256 0 -1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2375
timestamp 1644511149
transform 1 0 11408 0 -1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2376
timestamp 1644511149
transform 1 0 16560 0 -1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2377
timestamp 1644511149
transform 1 0 21712 0 -1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2378
timestamp 1644511149
transform 1 0 26864 0 -1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2379
timestamp 1644511149
transform 1 0 32016 0 -1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2380
timestamp 1644511149
transform 1 0 37168 0 -1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2381
timestamp 1644511149
transform 1 0 42320 0 -1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2382
timestamp 1644511149
transform 1 0 47472 0 -1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2383
timestamp 1644511149
transform 1 0 52624 0 -1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2384
timestamp 1644511149
transform 1 0 57776 0 -1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2385
timestamp 1644511149
transform 1 0 62928 0 -1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2386
timestamp 1644511149
transform 1 0 68080 0 -1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2387
timestamp 1644511149
transform 1 0 73232 0 -1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2388
timestamp 1644511149
transform 1 0 78384 0 -1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2389
timestamp 1644511149
transform 1 0 3680 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2390
timestamp 1644511149
transform 1 0 8832 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2391
timestamp 1644511149
transform 1 0 13984 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2392
timestamp 1644511149
transform 1 0 19136 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2393
timestamp 1644511149
transform 1 0 24288 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2394
timestamp 1644511149
transform 1 0 29440 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2395
timestamp 1644511149
transform 1 0 34592 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2396
timestamp 1644511149
transform 1 0 39744 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2397
timestamp 1644511149
transform 1 0 44896 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2398
timestamp 1644511149
transform 1 0 50048 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2399
timestamp 1644511149
transform 1 0 55200 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2400
timestamp 1644511149
transform 1 0 60352 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2401
timestamp 1644511149
transform 1 0 65504 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2402
timestamp 1644511149
transform 1 0 70656 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2403
timestamp 1644511149
transform 1 0 75808 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2404
timestamp 1644511149
transform 1 0 6256 0 -1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2405
timestamp 1644511149
transform 1 0 11408 0 -1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2406
timestamp 1644511149
transform 1 0 16560 0 -1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2407
timestamp 1644511149
transform 1 0 21712 0 -1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2408
timestamp 1644511149
transform 1 0 26864 0 -1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2409
timestamp 1644511149
transform 1 0 32016 0 -1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2410
timestamp 1644511149
transform 1 0 37168 0 -1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2411
timestamp 1644511149
transform 1 0 42320 0 -1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2412
timestamp 1644511149
transform 1 0 47472 0 -1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2413
timestamp 1644511149
transform 1 0 52624 0 -1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2414
timestamp 1644511149
transform 1 0 57776 0 -1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2415
timestamp 1644511149
transform 1 0 62928 0 -1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2416
timestamp 1644511149
transform 1 0 68080 0 -1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2417
timestamp 1644511149
transform 1 0 73232 0 -1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2418
timestamp 1644511149
transform 1 0 78384 0 -1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2419
timestamp 1644511149
transform 1 0 3680 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2420
timestamp 1644511149
transform 1 0 8832 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2421
timestamp 1644511149
transform 1 0 13984 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2422
timestamp 1644511149
transform 1 0 19136 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2423
timestamp 1644511149
transform 1 0 24288 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2424
timestamp 1644511149
transform 1 0 29440 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2425
timestamp 1644511149
transform 1 0 34592 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2426
timestamp 1644511149
transform 1 0 39744 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2427
timestamp 1644511149
transform 1 0 44896 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2428
timestamp 1644511149
transform 1 0 50048 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2429
timestamp 1644511149
transform 1 0 55200 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2430
timestamp 1644511149
transform 1 0 60352 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2431
timestamp 1644511149
transform 1 0 65504 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2432
timestamp 1644511149
transform 1 0 70656 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2433
timestamp 1644511149
transform 1 0 75808 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2434
timestamp 1644511149
transform 1 0 6256 0 -1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2435
timestamp 1644511149
transform 1 0 11408 0 -1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2436
timestamp 1644511149
transform 1 0 16560 0 -1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2437
timestamp 1644511149
transform 1 0 21712 0 -1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2438
timestamp 1644511149
transform 1 0 26864 0 -1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2439
timestamp 1644511149
transform 1 0 32016 0 -1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2440
timestamp 1644511149
transform 1 0 37168 0 -1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2441
timestamp 1644511149
transform 1 0 42320 0 -1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2442
timestamp 1644511149
transform 1 0 47472 0 -1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2443
timestamp 1644511149
transform 1 0 52624 0 -1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2444
timestamp 1644511149
transform 1 0 57776 0 -1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2445
timestamp 1644511149
transform 1 0 62928 0 -1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2446
timestamp 1644511149
transform 1 0 68080 0 -1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2447
timestamp 1644511149
transform 1 0 73232 0 -1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2448
timestamp 1644511149
transform 1 0 78384 0 -1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2449
timestamp 1644511149
transform 1 0 3680 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2450
timestamp 1644511149
transform 1 0 8832 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2451
timestamp 1644511149
transform 1 0 13984 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2452
timestamp 1644511149
transform 1 0 19136 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2453
timestamp 1644511149
transform 1 0 24288 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2454
timestamp 1644511149
transform 1 0 29440 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2455
timestamp 1644511149
transform 1 0 34592 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2456
timestamp 1644511149
transform 1 0 39744 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2457
timestamp 1644511149
transform 1 0 44896 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2458
timestamp 1644511149
transform 1 0 50048 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2459
timestamp 1644511149
transform 1 0 55200 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2460
timestamp 1644511149
transform 1 0 60352 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2461
timestamp 1644511149
transform 1 0 65504 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2462
timestamp 1644511149
transform 1 0 70656 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2463
timestamp 1644511149
transform 1 0 75808 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2464
timestamp 1644511149
transform 1 0 6256 0 -1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2465
timestamp 1644511149
transform 1 0 11408 0 -1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2466
timestamp 1644511149
transform 1 0 16560 0 -1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2467
timestamp 1644511149
transform 1 0 21712 0 -1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2468
timestamp 1644511149
transform 1 0 26864 0 -1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2469
timestamp 1644511149
transform 1 0 32016 0 -1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2470
timestamp 1644511149
transform 1 0 37168 0 -1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2471
timestamp 1644511149
transform 1 0 42320 0 -1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2472
timestamp 1644511149
transform 1 0 47472 0 -1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2473
timestamp 1644511149
transform 1 0 52624 0 -1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2474
timestamp 1644511149
transform 1 0 57776 0 -1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2475
timestamp 1644511149
transform 1 0 62928 0 -1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2476
timestamp 1644511149
transform 1 0 68080 0 -1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2477
timestamp 1644511149
transform 1 0 73232 0 -1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2478
timestamp 1644511149
transform 1 0 78384 0 -1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2479
timestamp 1644511149
transform 1 0 3680 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2480
timestamp 1644511149
transform 1 0 8832 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2481
timestamp 1644511149
transform 1 0 13984 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2482
timestamp 1644511149
transform 1 0 19136 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2483
timestamp 1644511149
transform 1 0 24288 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2484
timestamp 1644511149
transform 1 0 29440 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2485
timestamp 1644511149
transform 1 0 34592 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2486
timestamp 1644511149
transform 1 0 39744 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2487
timestamp 1644511149
transform 1 0 44896 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2488
timestamp 1644511149
transform 1 0 50048 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2489
timestamp 1644511149
transform 1 0 55200 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2490
timestamp 1644511149
transform 1 0 60352 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2491
timestamp 1644511149
transform 1 0 65504 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2492
timestamp 1644511149
transform 1 0 70656 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2493
timestamp 1644511149
transform 1 0 75808 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2494
timestamp 1644511149
transform 1 0 6256 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2495
timestamp 1644511149
transform 1 0 11408 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2496
timestamp 1644511149
transform 1 0 16560 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2497
timestamp 1644511149
transform 1 0 21712 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2498
timestamp 1644511149
transform 1 0 26864 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2499
timestamp 1644511149
transform 1 0 32016 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2500
timestamp 1644511149
transform 1 0 37168 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2501
timestamp 1644511149
transform 1 0 42320 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2502
timestamp 1644511149
transform 1 0 47472 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2503
timestamp 1644511149
transform 1 0 52624 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2504
timestamp 1644511149
transform 1 0 57776 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2505
timestamp 1644511149
transform 1 0 62928 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2506
timestamp 1644511149
transform 1 0 68080 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2507
timestamp 1644511149
transform 1 0 73232 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2508
timestamp 1644511149
transform 1 0 78384 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2509
timestamp 1644511149
transform 1 0 3680 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2510
timestamp 1644511149
transform 1 0 8832 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2511
timestamp 1644511149
transform 1 0 13984 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2512
timestamp 1644511149
transform 1 0 19136 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2513
timestamp 1644511149
transform 1 0 24288 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2514
timestamp 1644511149
transform 1 0 29440 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2515
timestamp 1644511149
transform 1 0 34592 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2516
timestamp 1644511149
transform 1 0 39744 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2517
timestamp 1644511149
transform 1 0 44896 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2518
timestamp 1644511149
transform 1 0 50048 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2519
timestamp 1644511149
transform 1 0 55200 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2520
timestamp 1644511149
transform 1 0 60352 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2521
timestamp 1644511149
transform 1 0 65504 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2522
timestamp 1644511149
transform 1 0 70656 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2523
timestamp 1644511149
transform 1 0 75808 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2524
timestamp 1644511149
transform 1 0 6256 0 -1 78336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2525
timestamp 1644511149
transform 1 0 11408 0 -1 78336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2526
timestamp 1644511149
transform 1 0 16560 0 -1 78336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2527
timestamp 1644511149
transform 1 0 21712 0 -1 78336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2528
timestamp 1644511149
transform 1 0 26864 0 -1 78336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2529
timestamp 1644511149
transform 1 0 32016 0 -1 78336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2530
timestamp 1644511149
transform 1 0 37168 0 -1 78336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2531
timestamp 1644511149
transform 1 0 42320 0 -1 78336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2532
timestamp 1644511149
transform 1 0 47472 0 -1 78336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2533
timestamp 1644511149
transform 1 0 52624 0 -1 78336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2534
timestamp 1644511149
transform 1 0 57776 0 -1 78336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2535
timestamp 1644511149
transform 1 0 62928 0 -1 78336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2536
timestamp 1644511149
transform 1 0 68080 0 -1 78336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2537
timestamp 1644511149
transform 1 0 73232 0 -1 78336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2538
timestamp 1644511149
transform 1 0 78384 0 -1 78336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2539
timestamp 1644511149
transform 1 0 3680 0 1 78336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2540
timestamp 1644511149
transform 1 0 8832 0 1 78336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2541
timestamp 1644511149
transform 1 0 13984 0 1 78336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2542
timestamp 1644511149
transform 1 0 19136 0 1 78336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2543
timestamp 1644511149
transform 1 0 24288 0 1 78336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2544
timestamp 1644511149
transform 1 0 29440 0 1 78336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2545
timestamp 1644511149
transform 1 0 34592 0 1 78336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2546
timestamp 1644511149
transform 1 0 39744 0 1 78336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2547
timestamp 1644511149
transform 1 0 44896 0 1 78336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2548
timestamp 1644511149
transform 1 0 50048 0 1 78336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2549
timestamp 1644511149
transform 1 0 55200 0 1 78336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2550
timestamp 1644511149
transform 1 0 60352 0 1 78336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2551
timestamp 1644511149
transform 1 0 65504 0 1 78336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2552
timestamp 1644511149
transform 1 0 70656 0 1 78336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2553
timestamp 1644511149
transform 1 0 75808 0 1 78336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2554
timestamp 1644511149
transform 1 0 6256 0 -1 79424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2555
timestamp 1644511149
transform 1 0 11408 0 -1 79424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2556
timestamp 1644511149
transform 1 0 16560 0 -1 79424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2557
timestamp 1644511149
transform 1 0 21712 0 -1 79424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2558
timestamp 1644511149
transform 1 0 26864 0 -1 79424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2559
timestamp 1644511149
transform 1 0 32016 0 -1 79424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2560
timestamp 1644511149
transform 1 0 37168 0 -1 79424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2561
timestamp 1644511149
transform 1 0 42320 0 -1 79424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2562
timestamp 1644511149
transform 1 0 47472 0 -1 79424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2563
timestamp 1644511149
transform 1 0 52624 0 -1 79424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2564
timestamp 1644511149
transform 1 0 57776 0 -1 79424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2565
timestamp 1644511149
transform 1 0 62928 0 -1 79424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2566
timestamp 1644511149
transform 1 0 68080 0 -1 79424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2567
timestamp 1644511149
transform 1 0 73232 0 -1 79424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2568
timestamp 1644511149
transform 1 0 78384 0 -1 79424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2569
timestamp 1644511149
transform 1 0 3680 0 1 79424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2570
timestamp 1644511149
transform 1 0 8832 0 1 79424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2571
timestamp 1644511149
transform 1 0 13984 0 1 79424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2572
timestamp 1644511149
transform 1 0 19136 0 1 79424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2573
timestamp 1644511149
transform 1 0 24288 0 1 79424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2574
timestamp 1644511149
transform 1 0 29440 0 1 79424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2575
timestamp 1644511149
transform 1 0 34592 0 1 79424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2576
timestamp 1644511149
transform 1 0 39744 0 1 79424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2577
timestamp 1644511149
transform 1 0 44896 0 1 79424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2578
timestamp 1644511149
transform 1 0 50048 0 1 79424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2579
timestamp 1644511149
transform 1 0 55200 0 1 79424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2580
timestamp 1644511149
transform 1 0 60352 0 1 79424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2581
timestamp 1644511149
transform 1 0 65504 0 1 79424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2582
timestamp 1644511149
transform 1 0 70656 0 1 79424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2583
timestamp 1644511149
transform 1 0 75808 0 1 79424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2584
timestamp 1644511149
transform 1 0 6256 0 -1 80512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2585
timestamp 1644511149
transform 1 0 11408 0 -1 80512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2586
timestamp 1644511149
transform 1 0 16560 0 -1 80512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2587
timestamp 1644511149
transform 1 0 21712 0 -1 80512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2588
timestamp 1644511149
transform 1 0 26864 0 -1 80512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2589
timestamp 1644511149
transform 1 0 32016 0 -1 80512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2590
timestamp 1644511149
transform 1 0 37168 0 -1 80512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2591
timestamp 1644511149
transform 1 0 42320 0 -1 80512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2592
timestamp 1644511149
transform 1 0 47472 0 -1 80512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2593
timestamp 1644511149
transform 1 0 52624 0 -1 80512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2594
timestamp 1644511149
transform 1 0 57776 0 -1 80512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2595
timestamp 1644511149
transform 1 0 62928 0 -1 80512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2596
timestamp 1644511149
transform 1 0 68080 0 -1 80512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2597
timestamp 1644511149
transform 1 0 73232 0 -1 80512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2598
timestamp 1644511149
transform 1 0 78384 0 -1 80512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2599
timestamp 1644511149
transform 1 0 3680 0 1 80512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2600
timestamp 1644511149
transform 1 0 8832 0 1 80512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2601
timestamp 1644511149
transform 1 0 13984 0 1 80512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2602
timestamp 1644511149
transform 1 0 19136 0 1 80512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2603
timestamp 1644511149
transform 1 0 24288 0 1 80512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2604
timestamp 1644511149
transform 1 0 29440 0 1 80512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2605
timestamp 1644511149
transform 1 0 34592 0 1 80512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2606
timestamp 1644511149
transform 1 0 39744 0 1 80512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2607
timestamp 1644511149
transform 1 0 44896 0 1 80512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2608
timestamp 1644511149
transform 1 0 50048 0 1 80512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2609
timestamp 1644511149
transform 1 0 55200 0 1 80512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2610
timestamp 1644511149
transform 1 0 60352 0 1 80512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2611
timestamp 1644511149
transform 1 0 65504 0 1 80512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2612
timestamp 1644511149
transform 1 0 70656 0 1 80512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2613
timestamp 1644511149
transform 1 0 75808 0 1 80512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2614
timestamp 1644511149
transform 1 0 6256 0 -1 81600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2615
timestamp 1644511149
transform 1 0 11408 0 -1 81600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2616
timestamp 1644511149
transform 1 0 16560 0 -1 81600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2617
timestamp 1644511149
transform 1 0 21712 0 -1 81600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2618
timestamp 1644511149
transform 1 0 26864 0 -1 81600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2619
timestamp 1644511149
transform 1 0 32016 0 -1 81600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2620
timestamp 1644511149
transform 1 0 37168 0 -1 81600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2621
timestamp 1644511149
transform 1 0 42320 0 -1 81600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2622
timestamp 1644511149
transform 1 0 47472 0 -1 81600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2623
timestamp 1644511149
transform 1 0 52624 0 -1 81600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2624
timestamp 1644511149
transform 1 0 57776 0 -1 81600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2625
timestamp 1644511149
transform 1 0 62928 0 -1 81600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2626
timestamp 1644511149
transform 1 0 68080 0 -1 81600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2627
timestamp 1644511149
transform 1 0 73232 0 -1 81600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2628
timestamp 1644511149
transform 1 0 78384 0 -1 81600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2629
timestamp 1644511149
transform 1 0 3680 0 1 81600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2630
timestamp 1644511149
transform 1 0 8832 0 1 81600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2631
timestamp 1644511149
transform 1 0 13984 0 1 81600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2632
timestamp 1644511149
transform 1 0 19136 0 1 81600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2633
timestamp 1644511149
transform 1 0 24288 0 1 81600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2634
timestamp 1644511149
transform 1 0 29440 0 1 81600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2635
timestamp 1644511149
transform 1 0 34592 0 1 81600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2636
timestamp 1644511149
transform 1 0 39744 0 1 81600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2637
timestamp 1644511149
transform 1 0 44896 0 1 81600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2638
timestamp 1644511149
transform 1 0 50048 0 1 81600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2639
timestamp 1644511149
transform 1 0 55200 0 1 81600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2640
timestamp 1644511149
transform 1 0 60352 0 1 81600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2641
timestamp 1644511149
transform 1 0 65504 0 1 81600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2642
timestamp 1644511149
transform 1 0 70656 0 1 81600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2643
timestamp 1644511149
transform 1 0 75808 0 1 81600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2644
timestamp 1644511149
transform 1 0 6256 0 -1 82688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2645
timestamp 1644511149
transform 1 0 11408 0 -1 82688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2646
timestamp 1644511149
transform 1 0 16560 0 -1 82688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2647
timestamp 1644511149
transform 1 0 21712 0 -1 82688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2648
timestamp 1644511149
transform 1 0 26864 0 -1 82688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2649
timestamp 1644511149
transform 1 0 32016 0 -1 82688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2650
timestamp 1644511149
transform 1 0 37168 0 -1 82688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2651
timestamp 1644511149
transform 1 0 42320 0 -1 82688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2652
timestamp 1644511149
transform 1 0 47472 0 -1 82688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2653
timestamp 1644511149
transform 1 0 52624 0 -1 82688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2654
timestamp 1644511149
transform 1 0 57776 0 -1 82688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2655
timestamp 1644511149
transform 1 0 62928 0 -1 82688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2656
timestamp 1644511149
transform 1 0 68080 0 -1 82688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2657
timestamp 1644511149
transform 1 0 73232 0 -1 82688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2658
timestamp 1644511149
transform 1 0 78384 0 -1 82688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2659
timestamp 1644511149
transform 1 0 3680 0 1 82688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2660
timestamp 1644511149
transform 1 0 8832 0 1 82688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2661
timestamp 1644511149
transform 1 0 13984 0 1 82688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2662
timestamp 1644511149
transform 1 0 19136 0 1 82688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2663
timestamp 1644511149
transform 1 0 24288 0 1 82688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2664
timestamp 1644511149
transform 1 0 29440 0 1 82688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2665
timestamp 1644511149
transform 1 0 34592 0 1 82688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2666
timestamp 1644511149
transform 1 0 39744 0 1 82688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2667
timestamp 1644511149
transform 1 0 44896 0 1 82688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2668
timestamp 1644511149
transform 1 0 50048 0 1 82688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2669
timestamp 1644511149
transform 1 0 55200 0 1 82688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2670
timestamp 1644511149
transform 1 0 60352 0 1 82688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2671
timestamp 1644511149
transform 1 0 65504 0 1 82688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2672
timestamp 1644511149
transform 1 0 70656 0 1 82688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2673
timestamp 1644511149
transform 1 0 75808 0 1 82688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2674
timestamp 1644511149
transform 1 0 6256 0 -1 83776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2675
timestamp 1644511149
transform 1 0 11408 0 -1 83776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2676
timestamp 1644511149
transform 1 0 16560 0 -1 83776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2677
timestamp 1644511149
transform 1 0 21712 0 -1 83776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2678
timestamp 1644511149
transform 1 0 26864 0 -1 83776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2679
timestamp 1644511149
transform 1 0 32016 0 -1 83776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2680
timestamp 1644511149
transform 1 0 37168 0 -1 83776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2681
timestamp 1644511149
transform 1 0 42320 0 -1 83776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2682
timestamp 1644511149
transform 1 0 47472 0 -1 83776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2683
timestamp 1644511149
transform 1 0 52624 0 -1 83776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2684
timestamp 1644511149
transform 1 0 57776 0 -1 83776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2685
timestamp 1644511149
transform 1 0 62928 0 -1 83776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2686
timestamp 1644511149
transform 1 0 68080 0 -1 83776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2687
timestamp 1644511149
transform 1 0 73232 0 -1 83776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2688
timestamp 1644511149
transform 1 0 78384 0 -1 83776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2689
timestamp 1644511149
transform 1 0 3680 0 1 83776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2690
timestamp 1644511149
transform 1 0 8832 0 1 83776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2691
timestamp 1644511149
transform 1 0 13984 0 1 83776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2692
timestamp 1644511149
transform 1 0 19136 0 1 83776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2693
timestamp 1644511149
transform 1 0 24288 0 1 83776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2694
timestamp 1644511149
transform 1 0 29440 0 1 83776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2695
timestamp 1644511149
transform 1 0 34592 0 1 83776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2696
timestamp 1644511149
transform 1 0 39744 0 1 83776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2697
timestamp 1644511149
transform 1 0 44896 0 1 83776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2698
timestamp 1644511149
transform 1 0 50048 0 1 83776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2699
timestamp 1644511149
transform 1 0 55200 0 1 83776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2700
timestamp 1644511149
transform 1 0 60352 0 1 83776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2701
timestamp 1644511149
transform 1 0 65504 0 1 83776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2702
timestamp 1644511149
transform 1 0 70656 0 1 83776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2703
timestamp 1644511149
transform 1 0 75808 0 1 83776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2704
timestamp 1644511149
transform 1 0 6256 0 -1 84864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2705
timestamp 1644511149
transform 1 0 11408 0 -1 84864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2706
timestamp 1644511149
transform 1 0 16560 0 -1 84864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2707
timestamp 1644511149
transform 1 0 21712 0 -1 84864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2708
timestamp 1644511149
transform 1 0 26864 0 -1 84864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2709
timestamp 1644511149
transform 1 0 32016 0 -1 84864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2710
timestamp 1644511149
transform 1 0 37168 0 -1 84864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2711
timestamp 1644511149
transform 1 0 42320 0 -1 84864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2712
timestamp 1644511149
transform 1 0 47472 0 -1 84864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2713
timestamp 1644511149
transform 1 0 52624 0 -1 84864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2714
timestamp 1644511149
transform 1 0 57776 0 -1 84864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2715
timestamp 1644511149
transform 1 0 62928 0 -1 84864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2716
timestamp 1644511149
transform 1 0 68080 0 -1 84864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2717
timestamp 1644511149
transform 1 0 73232 0 -1 84864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2718
timestamp 1644511149
transform 1 0 78384 0 -1 84864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2719
timestamp 1644511149
transform 1 0 3680 0 1 84864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2720
timestamp 1644511149
transform 1 0 8832 0 1 84864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2721
timestamp 1644511149
transform 1 0 13984 0 1 84864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2722
timestamp 1644511149
transform 1 0 19136 0 1 84864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2723
timestamp 1644511149
transform 1 0 24288 0 1 84864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2724
timestamp 1644511149
transform 1 0 29440 0 1 84864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2725
timestamp 1644511149
transform 1 0 34592 0 1 84864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2726
timestamp 1644511149
transform 1 0 39744 0 1 84864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2727
timestamp 1644511149
transform 1 0 44896 0 1 84864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2728
timestamp 1644511149
transform 1 0 50048 0 1 84864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2729
timestamp 1644511149
transform 1 0 55200 0 1 84864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2730
timestamp 1644511149
transform 1 0 60352 0 1 84864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2731
timestamp 1644511149
transform 1 0 65504 0 1 84864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2732
timestamp 1644511149
transform 1 0 70656 0 1 84864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2733
timestamp 1644511149
transform 1 0 75808 0 1 84864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2734
timestamp 1644511149
transform 1 0 6256 0 -1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2735
timestamp 1644511149
transform 1 0 11408 0 -1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2736
timestamp 1644511149
transform 1 0 16560 0 -1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2737
timestamp 1644511149
transform 1 0 21712 0 -1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2738
timestamp 1644511149
transform 1 0 26864 0 -1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2739
timestamp 1644511149
transform 1 0 32016 0 -1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2740
timestamp 1644511149
transform 1 0 37168 0 -1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2741
timestamp 1644511149
transform 1 0 42320 0 -1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2742
timestamp 1644511149
transform 1 0 47472 0 -1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2743
timestamp 1644511149
transform 1 0 52624 0 -1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2744
timestamp 1644511149
transform 1 0 57776 0 -1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2745
timestamp 1644511149
transform 1 0 62928 0 -1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2746
timestamp 1644511149
transform 1 0 68080 0 -1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2747
timestamp 1644511149
transform 1 0 73232 0 -1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2748
timestamp 1644511149
transform 1 0 78384 0 -1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2749
timestamp 1644511149
transform 1 0 3680 0 1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2750
timestamp 1644511149
transform 1 0 8832 0 1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2751
timestamp 1644511149
transform 1 0 13984 0 1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2752
timestamp 1644511149
transform 1 0 19136 0 1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2753
timestamp 1644511149
transform 1 0 24288 0 1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2754
timestamp 1644511149
transform 1 0 29440 0 1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2755
timestamp 1644511149
transform 1 0 34592 0 1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2756
timestamp 1644511149
transform 1 0 39744 0 1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2757
timestamp 1644511149
transform 1 0 44896 0 1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2758
timestamp 1644511149
transform 1 0 50048 0 1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2759
timestamp 1644511149
transform 1 0 55200 0 1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2760
timestamp 1644511149
transform 1 0 60352 0 1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2761
timestamp 1644511149
transform 1 0 65504 0 1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2762
timestamp 1644511149
transform 1 0 70656 0 1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2763
timestamp 1644511149
transform 1 0 75808 0 1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2764
timestamp 1644511149
transform 1 0 6256 0 -1 87040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2765
timestamp 1644511149
transform 1 0 11408 0 -1 87040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2766
timestamp 1644511149
transform 1 0 16560 0 -1 87040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2767
timestamp 1644511149
transform 1 0 21712 0 -1 87040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2768
timestamp 1644511149
transform 1 0 26864 0 -1 87040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2769
timestamp 1644511149
transform 1 0 32016 0 -1 87040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2770
timestamp 1644511149
transform 1 0 37168 0 -1 87040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2771
timestamp 1644511149
transform 1 0 42320 0 -1 87040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2772
timestamp 1644511149
transform 1 0 47472 0 -1 87040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2773
timestamp 1644511149
transform 1 0 52624 0 -1 87040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2774
timestamp 1644511149
transform 1 0 57776 0 -1 87040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2775
timestamp 1644511149
transform 1 0 62928 0 -1 87040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2776
timestamp 1644511149
transform 1 0 68080 0 -1 87040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2777
timestamp 1644511149
transform 1 0 73232 0 -1 87040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2778
timestamp 1644511149
transform 1 0 78384 0 -1 87040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2779
timestamp 1644511149
transform 1 0 3680 0 1 87040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2780
timestamp 1644511149
transform 1 0 8832 0 1 87040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2781
timestamp 1644511149
transform 1 0 13984 0 1 87040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2782
timestamp 1644511149
transform 1 0 19136 0 1 87040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2783
timestamp 1644511149
transform 1 0 24288 0 1 87040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2784
timestamp 1644511149
transform 1 0 29440 0 1 87040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2785
timestamp 1644511149
transform 1 0 34592 0 1 87040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2786
timestamp 1644511149
transform 1 0 39744 0 1 87040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2787
timestamp 1644511149
transform 1 0 44896 0 1 87040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2788
timestamp 1644511149
transform 1 0 50048 0 1 87040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2789
timestamp 1644511149
transform 1 0 55200 0 1 87040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2790
timestamp 1644511149
transform 1 0 60352 0 1 87040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2791
timestamp 1644511149
transform 1 0 65504 0 1 87040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2792
timestamp 1644511149
transform 1 0 70656 0 1 87040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2793
timestamp 1644511149
transform 1 0 75808 0 1 87040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2794
timestamp 1644511149
transform 1 0 6256 0 -1 88128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2795
timestamp 1644511149
transform 1 0 11408 0 -1 88128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2796
timestamp 1644511149
transform 1 0 16560 0 -1 88128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2797
timestamp 1644511149
transform 1 0 21712 0 -1 88128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2798
timestamp 1644511149
transform 1 0 26864 0 -1 88128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2799
timestamp 1644511149
transform 1 0 32016 0 -1 88128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2800
timestamp 1644511149
transform 1 0 37168 0 -1 88128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2801
timestamp 1644511149
transform 1 0 42320 0 -1 88128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2802
timestamp 1644511149
transform 1 0 47472 0 -1 88128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2803
timestamp 1644511149
transform 1 0 52624 0 -1 88128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2804
timestamp 1644511149
transform 1 0 57776 0 -1 88128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2805
timestamp 1644511149
transform 1 0 62928 0 -1 88128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2806
timestamp 1644511149
transform 1 0 68080 0 -1 88128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2807
timestamp 1644511149
transform 1 0 73232 0 -1 88128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2808
timestamp 1644511149
transform 1 0 78384 0 -1 88128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2809
timestamp 1644511149
transform 1 0 3680 0 1 88128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2810
timestamp 1644511149
transform 1 0 8832 0 1 88128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2811
timestamp 1644511149
transform 1 0 13984 0 1 88128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2812
timestamp 1644511149
transform 1 0 19136 0 1 88128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2813
timestamp 1644511149
transform 1 0 24288 0 1 88128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2814
timestamp 1644511149
transform 1 0 29440 0 1 88128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2815
timestamp 1644511149
transform 1 0 34592 0 1 88128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2816
timestamp 1644511149
transform 1 0 39744 0 1 88128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2817
timestamp 1644511149
transform 1 0 44896 0 1 88128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2818
timestamp 1644511149
transform 1 0 50048 0 1 88128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2819
timestamp 1644511149
transform 1 0 55200 0 1 88128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2820
timestamp 1644511149
transform 1 0 60352 0 1 88128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2821
timestamp 1644511149
transform 1 0 65504 0 1 88128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2822
timestamp 1644511149
transform 1 0 70656 0 1 88128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2823
timestamp 1644511149
transform 1 0 75808 0 1 88128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2824
timestamp 1644511149
transform 1 0 6256 0 -1 89216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2825
timestamp 1644511149
transform 1 0 11408 0 -1 89216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2826
timestamp 1644511149
transform 1 0 16560 0 -1 89216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2827
timestamp 1644511149
transform 1 0 21712 0 -1 89216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2828
timestamp 1644511149
transform 1 0 26864 0 -1 89216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2829
timestamp 1644511149
transform 1 0 32016 0 -1 89216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2830
timestamp 1644511149
transform 1 0 37168 0 -1 89216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2831
timestamp 1644511149
transform 1 0 42320 0 -1 89216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2832
timestamp 1644511149
transform 1 0 47472 0 -1 89216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2833
timestamp 1644511149
transform 1 0 52624 0 -1 89216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2834
timestamp 1644511149
transform 1 0 57776 0 -1 89216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2835
timestamp 1644511149
transform 1 0 62928 0 -1 89216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2836
timestamp 1644511149
transform 1 0 68080 0 -1 89216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2837
timestamp 1644511149
transform 1 0 73232 0 -1 89216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2838
timestamp 1644511149
transform 1 0 78384 0 -1 89216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2839
timestamp 1644511149
transform 1 0 3680 0 1 89216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2840
timestamp 1644511149
transform 1 0 8832 0 1 89216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2841
timestamp 1644511149
transform 1 0 13984 0 1 89216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2842
timestamp 1644511149
transform 1 0 19136 0 1 89216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2843
timestamp 1644511149
transform 1 0 24288 0 1 89216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2844
timestamp 1644511149
transform 1 0 29440 0 1 89216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2845
timestamp 1644511149
transform 1 0 34592 0 1 89216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2846
timestamp 1644511149
transform 1 0 39744 0 1 89216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2847
timestamp 1644511149
transform 1 0 44896 0 1 89216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2848
timestamp 1644511149
transform 1 0 50048 0 1 89216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2849
timestamp 1644511149
transform 1 0 55200 0 1 89216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2850
timestamp 1644511149
transform 1 0 60352 0 1 89216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2851
timestamp 1644511149
transform 1 0 65504 0 1 89216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2852
timestamp 1644511149
transform 1 0 70656 0 1 89216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2853
timestamp 1644511149
transform 1 0 75808 0 1 89216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2854
timestamp 1644511149
transform 1 0 6256 0 -1 90304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2855
timestamp 1644511149
transform 1 0 11408 0 -1 90304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2856
timestamp 1644511149
transform 1 0 16560 0 -1 90304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2857
timestamp 1644511149
transform 1 0 21712 0 -1 90304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2858
timestamp 1644511149
transform 1 0 26864 0 -1 90304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2859
timestamp 1644511149
transform 1 0 32016 0 -1 90304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2860
timestamp 1644511149
transform 1 0 37168 0 -1 90304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2861
timestamp 1644511149
transform 1 0 42320 0 -1 90304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2862
timestamp 1644511149
transform 1 0 47472 0 -1 90304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2863
timestamp 1644511149
transform 1 0 52624 0 -1 90304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2864
timestamp 1644511149
transform 1 0 57776 0 -1 90304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2865
timestamp 1644511149
transform 1 0 62928 0 -1 90304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2866
timestamp 1644511149
transform 1 0 68080 0 -1 90304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2867
timestamp 1644511149
transform 1 0 73232 0 -1 90304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2868
timestamp 1644511149
transform 1 0 78384 0 -1 90304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2869
timestamp 1644511149
transform 1 0 3680 0 1 90304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2870
timestamp 1644511149
transform 1 0 8832 0 1 90304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2871
timestamp 1644511149
transform 1 0 13984 0 1 90304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2872
timestamp 1644511149
transform 1 0 19136 0 1 90304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2873
timestamp 1644511149
transform 1 0 24288 0 1 90304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2874
timestamp 1644511149
transform 1 0 29440 0 1 90304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2875
timestamp 1644511149
transform 1 0 34592 0 1 90304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2876
timestamp 1644511149
transform 1 0 39744 0 1 90304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2877
timestamp 1644511149
transform 1 0 44896 0 1 90304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2878
timestamp 1644511149
transform 1 0 50048 0 1 90304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2879
timestamp 1644511149
transform 1 0 55200 0 1 90304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2880
timestamp 1644511149
transform 1 0 60352 0 1 90304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2881
timestamp 1644511149
transform 1 0 65504 0 1 90304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2882
timestamp 1644511149
transform 1 0 70656 0 1 90304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2883
timestamp 1644511149
transform 1 0 75808 0 1 90304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2884
timestamp 1644511149
transform 1 0 6256 0 -1 91392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2885
timestamp 1644511149
transform 1 0 11408 0 -1 91392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2886
timestamp 1644511149
transform 1 0 16560 0 -1 91392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2887
timestamp 1644511149
transform 1 0 21712 0 -1 91392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2888
timestamp 1644511149
transform 1 0 26864 0 -1 91392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2889
timestamp 1644511149
transform 1 0 32016 0 -1 91392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2890
timestamp 1644511149
transform 1 0 37168 0 -1 91392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2891
timestamp 1644511149
transform 1 0 42320 0 -1 91392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2892
timestamp 1644511149
transform 1 0 47472 0 -1 91392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2893
timestamp 1644511149
transform 1 0 52624 0 -1 91392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2894
timestamp 1644511149
transform 1 0 57776 0 -1 91392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2895
timestamp 1644511149
transform 1 0 62928 0 -1 91392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2896
timestamp 1644511149
transform 1 0 68080 0 -1 91392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2897
timestamp 1644511149
transform 1 0 73232 0 -1 91392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2898
timestamp 1644511149
transform 1 0 78384 0 -1 91392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2899
timestamp 1644511149
transform 1 0 3680 0 1 91392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2900
timestamp 1644511149
transform 1 0 8832 0 1 91392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2901
timestamp 1644511149
transform 1 0 13984 0 1 91392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2902
timestamp 1644511149
transform 1 0 19136 0 1 91392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2903
timestamp 1644511149
transform 1 0 24288 0 1 91392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2904
timestamp 1644511149
transform 1 0 29440 0 1 91392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2905
timestamp 1644511149
transform 1 0 34592 0 1 91392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2906
timestamp 1644511149
transform 1 0 39744 0 1 91392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2907
timestamp 1644511149
transform 1 0 44896 0 1 91392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2908
timestamp 1644511149
transform 1 0 50048 0 1 91392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2909
timestamp 1644511149
transform 1 0 55200 0 1 91392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2910
timestamp 1644511149
transform 1 0 60352 0 1 91392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2911
timestamp 1644511149
transform 1 0 65504 0 1 91392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2912
timestamp 1644511149
transform 1 0 70656 0 1 91392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2913
timestamp 1644511149
transform 1 0 75808 0 1 91392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2914
timestamp 1644511149
transform 1 0 6256 0 -1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2915
timestamp 1644511149
transform 1 0 11408 0 -1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2916
timestamp 1644511149
transform 1 0 16560 0 -1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2917
timestamp 1644511149
transform 1 0 21712 0 -1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2918
timestamp 1644511149
transform 1 0 26864 0 -1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2919
timestamp 1644511149
transform 1 0 32016 0 -1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2920
timestamp 1644511149
transform 1 0 37168 0 -1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2921
timestamp 1644511149
transform 1 0 42320 0 -1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2922
timestamp 1644511149
transform 1 0 47472 0 -1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2923
timestamp 1644511149
transform 1 0 52624 0 -1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2924
timestamp 1644511149
transform 1 0 57776 0 -1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2925
timestamp 1644511149
transform 1 0 62928 0 -1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2926
timestamp 1644511149
transform 1 0 68080 0 -1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2927
timestamp 1644511149
transform 1 0 73232 0 -1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2928
timestamp 1644511149
transform 1 0 78384 0 -1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2929
timestamp 1644511149
transform 1 0 3680 0 1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2930
timestamp 1644511149
transform 1 0 8832 0 1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2931
timestamp 1644511149
transform 1 0 13984 0 1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2932
timestamp 1644511149
transform 1 0 19136 0 1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2933
timestamp 1644511149
transform 1 0 24288 0 1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2934
timestamp 1644511149
transform 1 0 29440 0 1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2935
timestamp 1644511149
transform 1 0 34592 0 1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2936
timestamp 1644511149
transform 1 0 39744 0 1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2937
timestamp 1644511149
transform 1 0 44896 0 1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2938
timestamp 1644511149
transform 1 0 50048 0 1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2939
timestamp 1644511149
transform 1 0 55200 0 1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2940
timestamp 1644511149
transform 1 0 60352 0 1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2941
timestamp 1644511149
transform 1 0 65504 0 1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2942
timestamp 1644511149
transform 1 0 70656 0 1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2943
timestamp 1644511149
transform 1 0 75808 0 1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2944
timestamp 1644511149
transform 1 0 6256 0 -1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2945
timestamp 1644511149
transform 1 0 11408 0 -1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2946
timestamp 1644511149
transform 1 0 16560 0 -1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2947
timestamp 1644511149
transform 1 0 21712 0 -1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2948
timestamp 1644511149
transform 1 0 26864 0 -1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2949
timestamp 1644511149
transform 1 0 32016 0 -1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2950
timestamp 1644511149
transform 1 0 37168 0 -1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2951
timestamp 1644511149
transform 1 0 42320 0 -1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2952
timestamp 1644511149
transform 1 0 47472 0 -1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2953
timestamp 1644511149
transform 1 0 52624 0 -1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2954
timestamp 1644511149
transform 1 0 57776 0 -1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2955
timestamp 1644511149
transform 1 0 62928 0 -1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2956
timestamp 1644511149
transform 1 0 68080 0 -1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2957
timestamp 1644511149
transform 1 0 73232 0 -1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2958
timestamp 1644511149
transform 1 0 78384 0 -1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2959
timestamp 1644511149
transform 1 0 3680 0 1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2960
timestamp 1644511149
transform 1 0 8832 0 1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2961
timestamp 1644511149
transform 1 0 13984 0 1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2962
timestamp 1644511149
transform 1 0 19136 0 1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2963
timestamp 1644511149
transform 1 0 24288 0 1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2964
timestamp 1644511149
transform 1 0 29440 0 1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2965
timestamp 1644511149
transform 1 0 34592 0 1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2966
timestamp 1644511149
transform 1 0 39744 0 1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2967
timestamp 1644511149
transform 1 0 44896 0 1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2968
timestamp 1644511149
transform 1 0 50048 0 1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2969
timestamp 1644511149
transform 1 0 55200 0 1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2970
timestamp 1644511149
transform 1 0 60352 0 1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2971
timestamp 1644511149
transform 1 0 65504 0 1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2972
timestamp 1644511149
transform 1 0 70656 0 1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2973
timestamp 1644511149
transform 1 0 75808 0 1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2974
timestamp 1644511149
transform 1 0 6256 0 -1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2975
timestamp 1644511149
transform 1 0 11408 0 -1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2976
timestamp 1644511149
transform 1 0 16560 0 -1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2977
timestamp 1644511149
transform 1 0 21712 0 -1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2978
timestamp 1644511149
transform 1 0 26864 0 -1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2979
timestamp 1644511149
transform 1 0 32016 0 -1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2980
timestamp 1644511149
transform 1 0 37168 0 -1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2981
timestamp 1644511149
transform 1 0 42320 0 -1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2982
timestamp 1644511149
transform 1 0 47472 0 -1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2983
timestamp 1644511149
transform 1 0 52624 0 -1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2984
timestamp 1644511149
transform 1 0 57776 0 -1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2985
timestamp 1644511149
transform 1 0 62928 0 -1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2986
timestamp 1644511149
transform 1 0 68080 0 -1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2987
timestamp 1644511149
transform 1 0 73232 0 -1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2988
timestamp 1644511149
transform 1 0 78384 0 -1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2989
timestamp 1644511149
transform 1 0 3680 0 1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2990
timestamp 1644511149
transform 1 0 8832 0 1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2991
timestamp 1644511149
transform 1 0 13984 0 1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2992
timestamp 1644511149
transform 1 0 19136 0 1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2993
timestamp 1644511149
transform 1 0 24288 0 1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2994
timestamp 1644511149
transform 1 0 29440 0 1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2995
timestamp 1644511149
transform 1 0 34592 0 1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2996
timestamp 1644511149
transform 1 0 39744 0 1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2997
timestamp 1644511149
transform 1 0 44896 0 1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2998
timestamp 1644511149
transform 1 0 50048 0 1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2999
timestamp 1644511149
transform 1 0 55200 0 1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3000
timestamp 1644511149
transform 1 0 60352 0 1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3001
timestamp 1644511149
transform 1 0 65504 0 1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3002
timestamp 1644511149
transform 1 0 70656 0 1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3003
timestamp 1644511149
transform 1 0 75808 0 1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3004
timestamp 1644511149
transform 1 0 6256 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3005
timestamp 1644511149
transform 1 0 11408 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3006
timestamp 1644511149
transform 1 0 16560 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3007
timestamp 1644511149
transform 1 0 21712 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3008
timestamp 1644511149
transform 1 0 26864 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3009
timestamp 1644511149
transform 1 0 32016 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3010
timestamp 1644511149
transform 1 0 37168 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3011
timestamp 1644511149
transform 1 0 42320 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3012
timestamp 1644511149
transform 1 0 47472 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3013
timestamp 1644511149
transform 1 0 52624 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3014
timestamp 1644511149
transform 1 0 57776 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3015
timestamp 1644511149
transform 1 0 62928 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3016
timestamp 1644511149
transform 1 0 68080 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3017
timestamp 1644511149
transform 1 0 73232 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3018
timestamp 1644511149
transform 1 0 78384 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3019
timestamp 1644511149
transform 1 0 3680 0 1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3020
timestamp 1644511149
transform 1 0 8832 0 1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3021
timestamp 1644511149
transform 1 0 13984 0 1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3022
timestamp 1644511149
transform 1 0 19136 0 1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3023
timestamp 1644511149
transform 1 0 24288 0 1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3024
timestamp 1644511149
transform 1 0 29440 0 1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3025
timestamp 1644511149
transform 1 0 34592 0 1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3026
timestamp 1644511149
transform 1 0 39744 0 1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3027
timestamp 1644511149
transform 1 0 44896 0 1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3028
timestamp 1644511149
transform 1 0 50048 0 1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3029
timestamp 1644511149
transform 1 0 55200 0 1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3030
timestamp 1644511149
transform 1 0 60352 0 1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3031
timestamp 1644511149
transform 1 0 65504 0 1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3032
timestamp 1644511149
transform 1 0 70656 0 1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3033
timestamp 1644511149
transform 1 0 75808 0 1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3034
timestamp 1644511149
transform 1 0 6256 0 -1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3035
timestamp 1644511149
transform 1 0 11408 0 -1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3036
timestamp 1644511149
transform 1 0 16560 0 -1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3037
timestamp 1644511149
transform 1 0 21712 0 -1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3038
timestamp 1644511149
transform 1 0 26864 0 -1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3039
timestamp 1644511149
transform 1 0 32016 0 -1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3040
timestamp 1644511149
transform 1 0 37168 0 -1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3041
timestamp 1644511149
transform 1 0 42320 0 -1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3042
timestamp 1644511149
transform 1 0 47472 0 -1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3043
timestamp 1644511149
transform 1 0 52624 0 -1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3044
timestamp 1644511149
transform 1 0 57776 0 -1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3045
timestamp 1644511149
transform 1 0 62928 0 -1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3046
timestamp 1644511149
transform 1 0 68080 0 -1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3047
timestamp 1644511149
transform 1 0 73232 0 -1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3048
timestamp 1644511149
transform 1 0 78384 0 -1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3049
timestamp 1644511149
transform 1 0 3680 0 1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3050
timestamp 1644511149
transform 1 0 8832 0 1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3051
timestamp 1644511149
transform 1 0 13984 0 1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3052
timestamp 1644511149
transform 1 0 19136 0 1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3053
timestamp 1644511149
transform 1 0 24288 0 1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3054
timestamp 1644511149
transform 1 0 29440 0 1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3055
timestamp 1644511149
transform 1 0 34592 0 1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3056
timestamp 1644511149
transform 1 0 39744 0 1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3057
timestamp 1644511149
transform 1 0 44896 0 1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3058
timestamp 1644511149
transform 1 0 50048 0 1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3059
timestamp 1644511149
transform 1 0 55200 0 1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3060
timestamp 1644511149
transform 1 0 60352 0 1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3061
timestamp 1644511149
transform 1 0 65504 0 1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3062
timestamp 1644511149
transform 1 0 70656 0 1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3063
timestamp 1644511149
transform 1 0 75808 0 1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3064
timestamp 1644511149
transform 1 0 6256 0 -1 97920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3065
timestamp 1644511149
transform 1 0 11408 0 -1 97920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3066
timestamp 1644511149
transform 1 0 16560 0 -1 97920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3067
timestamp 1644511149
transform 1 0 21712 0 -1 97920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3068
timestamp 1644511149
transform 1 0 26864 0 -1 97920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3069
timestamp 1644511149
transform 1 0 32016 0 -1 97920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3070
timestamp 1644511149
transform 1 0 37168 0 -1 97920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3071
timestamp 1644511149
transform 1 0 42320 0 -1 97920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3072
timestamp 1644511149
transform 1 0 47472 0 -1 97920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3073
timestamp 1644511149
transform 1 0 52624 0 -1 97920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3074
timestamp 1644511149
transform 1 0 57776 0 -1 97920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3075
timestamp 1644511149
transform 1 0 62928 0 -1 97920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3076
timestamp 1644511149
transform 1 0 68080 0 -1 97920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3077
timestamp 1644511149
transform 1 0 73232 0 -1 97920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3078
timestamp 1644511149
transform 1 0 78384 0 -1 97920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3079
timestamp 1644511149
transform 1 0 3680 0 1 97920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3080
timestamp 1644511149
transform 1 0 8832 0 1 97920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3081
timestamp 1644511149
transform 1 0 13984 0 1 97920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3082
timestamp 1644511149
transform 1 0 19136 0 1 97920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3083
timestamp 1644511149
transform 1 0 24288 0 1 97920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3084
timestamp 1644511149
transform 1 0 29440 0 1 97920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3085
timestamp 1644511149
transform 1 0 34592 0 1 97920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3086
timestamp 1644511149
transform 1 0 39744 0 1 97920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3087
timestamp 1644511149
transform 1 0 44896 0 1 97920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3088
timestamp 1644511149
transform 1 0 50048 0 1 97920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3089
timestamp 1644511149
transform 1 0 55200 0 1 97920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3090
timestamp 1644511149
transform 1 0 60352 0 1 97920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3091
timestamp 1644511149
transform 1 0 65504 0 1 97920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3092
timestamp 1644511149
transform 1 0 70656 0 1 97920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3093
timestamp 1644511149
transform 1 0 75808 0 1 97920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3094
timestamp 1644511149
transform 1 0 6256 0 -1 99008
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3095
timestamp 1644511149
transform 1 0 11408 0 -1 99008
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3096
timestamp 1644511149
transform 1 0 16560 0 -1 99008
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3097
timestamp 1644511149
transform 1 0 21712 0 -1 99008
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3098
timestamp 1644511149
transform 1 0 26864 0 -1 99008
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3099
timestamp 1644511149
transform 1 0 32016 0 -1 99008
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3100
timestamp 1644511149
transform 1 0 37168 0 -1 99008
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3101
timestamp 1644511149
transform 1 0 42320 0 -1 99008
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3102
timestamp 1644511149
transform 1 0 47472 0 -1 99008
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3103
timestamp 1644511149
transform 1 0 52624 0 -1 99008
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3104
timestamp 1644511149
transform 1 0 57776 0 -1 99008
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3105
timestamp 1644511149
transform 1 0 62928 0 -1 99008
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3106
timestamp 1644511149
transform 1 0 68080 0 -1 99008
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3107
timestamp 1644511149
transform 1 0 73232 0 -1 99008
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3108
timestamp 1644511149
transform 1 0 78384 0 -1 99008
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3109
timestamp 1644511149
transform 1 0 3680 0 1 99008
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3110
timestamp 1644511149
transform 1 0 8832 0 1 99008
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3111
timestamp 1644511149
transform 1 0 13984 0 1 99008
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3112
timestamp 1644511149
transform 1 0 19136 0 1 99008
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3113
timestamp 1644511149
transform 1 0 24288 0 1 99008
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3114
timestamp 1644511149
transform 1 0 29440 0 1 99008
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3115
timestamp 1644511149
transform 1 0 34592 0 1 99008
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3116
timestamp 1644511149
transform 1 0 39744 0 1 99008
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3117
timestamp 1644511149
transform 1 0 44896 0 1 99008
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3118
timestamp 1644511149
transform 1 0 50048 0 1 99008
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3119
timestamp 1644511149
transform 1 0 55200 0 1 99008
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3120
timestamp 1644511149
transform 1 0 60352 0 1 99008
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3121
timestamp 1644511149
transform 1 0 65504 0 1 99008
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3122
timestamp 1644511149
transform 1 0 70656 0 1 99008
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3123
timestamp 1644511149
transform 1 0 75808 0 1 99008
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3124
timestamp 1644511149
transform 1 0 6256 0 -1 100096
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3125
timestamp 1644511149
transform 1 0 11408 0 -1 100096
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3126
timestamp 1644511149
transform 1 0 16560 0 -1 100096
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3127
timestamp 1644511149
transform 1 0 21712 0 -1 100096
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3128
timestamp 1644511149
transform 1 0 26864 0 -1 100096
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3129
timestamp 1644511149
transform 1 0 32016 0 -1 100096
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3130
timestamp 1644511149
transform 1 0 37168 0 -1 100096
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3131
timestamp 1644511149
transform 1 0 42320 0 -1 100096
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3132
timestamp 1644511149
transform 1 0 47472 0 -1 100096
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3133
timestamp 1644511149
transform 1 0 52624 0 -1 100096
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3134
timestamp 1644511149
transform 1 0 57776 0 -1 100096
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3135
timestamp 1644511149
transform 1 0 62928 0 -1 100096
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3136
timestamp 1644511149
transform 1 0 68080 0 -1 100096
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3137
timestamp 1644511149
transform 1 0 73232 0 -1 100096
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3138
timestamp 1644511149
transform 1 0 78384 0 -1 100096
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3139
timestamp 1644511149
transform 1 0 3680 0 1 100096
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3140
timestamp 1644511149
transform 1 0 8832 0 1 100096
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3141
timestamp 1644511149
transform 1 0 13984 0 1 100096
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3142
timestamp 1644511149
transform 1 0 19136 0 1 100096
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3143
timestamp 1644511149
transform 1 0 24288 0 1 100096
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3144
timestamp 1644511149
transform 1 0 29440 0 1 100096
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3145
timestamp 1644511149
transform 1 0 34592 0 1 100096
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3146
timestamp 1644511149
transform 1 0 39744 0 1 100096
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3147
timestamp 1644511149
transform 1 0 44896 0 1 100096
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3148
timestamp 1644511149
transform 1 0 50048 0 1 100096
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3149
timestamp 1644511149
transform 1 0 55200 0 1 100096
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3150
timestamp 1644511149
transform 1 0 60352 0 1 100096
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3151
timestamp 1644511149
transform 1 0 65504 0 1 100096
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3152
timestamp 1644511149
transform 1 0 70656 0 1 100096
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3153
timestamp 1644511149
transform 1 0 75808 0 1 100096
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3154
timestamp 1644511149
transform 1 0 6256 0 -1 101184
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3155
timestamp 1644511149
transform 1 0 11408 0 -1 101184
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3156
timestamp 1644511149
transform 1 0 16560 0 -1 101184
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3157
timestamp 1644511149
transform 1 0 21712 0 -1 101184
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3158
timestamp 1644511149
transform 1 0 26864 0 -1 101184
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3159
timestamp 1644511149
transform 1 0 32016 0 -1 101184
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3160
timestamp 1644511149
transform 1 0 37168 0 -1 101184
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3161
timestamp 1644511149
transform 1 0 42320 0 -1 101184
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3162
timestamp 1644511149
transform 1 0 47472 0 -1 101184
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3163
timestamp 1644511149
transform 1 0 52624 0 -1 101184
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3164
timestamp 1644511149
transform 1 0 57776 0 -1 101184
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3165
timestamp 1644511149
transform 1 0 62928 0 -1 101184
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3166
timestamp 1644511149
transform 1 0 68080 0 -1 101184
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3167
timestamp 1644511149
transform 1 0 73232 0 -1 101184
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3168
timestamp 1644511149
transform 1 0 78384 0 -1 101184
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3169
timestamp 1644511149
transform 1 0 3680 0 1 101184
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3170
timestamp 1644511149
transform 1 0 8832 0 1 101184
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3171
timestamp 1644511149
transform 1 0 13984 0 1 101184
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3172
timestamp 1644511149
transform 1 0 19136 0 1 101184
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3173
timestamp 1644511149
transform 1 0 24288 0 1 101184
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3174
timestamp 1644511149
transform 1 0 29440 0 1 101184
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3175
timestamp 1644511149
transform 1 0 34592 0 1 101184
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3176
timestamp 1644511149
transform 1 0 39744 0 1 101184
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3177
timestamp 1644511149
transform 1 0 44896 0 1 101184
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3178
timestamp 1644511149
transform 1 0 50048 0 1 101184
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3179
timestamp 1644511149
transform 1 0 55200 0 1 101184
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3180
timestamp 1644511149
transform 1 0 60352 0 1 101184
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3181
timestamp 1644511149
transform 1 0 65504 0 1 101184
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3182
timestamp 1644511149
transform 1 0 70656 0 1 101184
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3183
timestamp 1644511149
transform 1 0 75808 0 1 101184
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3184
timestamp 1644511149
transform 1 0 6256 0 -1 102272
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3185
timestamp 1644511149
transform 1 0 11408 0 -1 102272
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3186
timestamp 1644511149
transform 1 0 16560 0 -1 102272
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3187
timestamp 1644511149
transform 1 0 21712 0 -1 102272
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3188
timestamp 1644511149
transform 1 0 26864 0 -1 102272
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3189
timestamp 1644511149
transform 1 0 32016 0 -1 102272
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3190
timestamp 1644511149
transform 1 0 37168 0 -1 102272
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3191
timestamp 1644511149
transform 1 0 42320 0 -1 102272
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3192
timestamp 1644511149
transform 1 0 47472 0 -1 102272
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3193
timestamp 1644511149
transform 1 0 52624 0 -1 102272
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3194
timestamp 1644511149
transform 1 0 57776 0 -1 102272
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3195
timestamp 1644511149
transform 1 0 62928 0 -1 102272
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3196
timestamp 1644511149
transform 1 0 68080 0 -1 102272
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3197
timestamp 1644511149
transform 1 0 73232 0 -1 102272
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3198
timestamp 1644511149
transform 1 0 78384 0 -1 102272
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3199
timestamp 1644511149
transform 1 0 3680 0 1 102272
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3200
timestamp 1644511149
transform 1 0 8832 0 1 102272
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3201
timestamp 1644511149
transform 1 0 13984 0 1 102272
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3202
timestamp 1644511149
transform 1 0 19136 0 1 102272
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3203
timestamp 1644511149
transform 1 0 24288 0 1 102272
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3204
timestamp 1644511149
transform 1 0 29440 0 1 102272
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3205
timestamp 1644511149
transform 1 0 34592 0 1 102272
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3206
timestamp 1644511149
transform 1 0 39744 0 1 102272
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3207
timestamp 1644511149
transform 1 0 44896 0 1 102272
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3208
timestamp 1644511149
transform 1 0 50048 0 1 102272
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3209
timestamp 1644511149
transform 1 0 55200 0 1 102272
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3210
timestamp 1644511149
transform 1 0 60352 0 1 102272
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3211
timestamp 1644511149
transform 1 0 65504 0 1 102272
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3212
timestamp 1644511149
transform 1 0 70656 0 1 102272
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3213
timestamp 1644511149
transform 1 0 75808 0 1 102272
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3214
timestamp 1644511149
transform 1 0 6256 0 -1 103360
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3215
timestamp 1644511149
transform 1 0 11408 0 -1 103360
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3216
timestamp 1644511149
transform 1 0 16560 0 -1 103360
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3217
timestamp 1644511149
transform 1 0 21712 0 -1 103360
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3218
timestamp 1644511149
transform 1 0 26864 0 -1 103360
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3219
timestamp 1644511149
transform 1 0 32016 0 -1 103360
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3220
timestamp 1644511149
transform 1 0 37168 0 -1 103360
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3221
timestamp 1644511149
transform 1 0 42320 0 -1 103360
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3222
timestamp 1644511149
transform 1 0 47472 0 -1 103360
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3223
timestamp 1644511149
transform 1 0 52624 0 -1 103360
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3224
timestamp 1644511149
transform 1 0 57776 0 -1 103360
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3225
timestamp 1644511149
transform 1 0 62928 0 -1 103360
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3226
timestamp 1644511149
transform 1 0 68080 0 -1 103360
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3227
timestamp 1644511149
transform 1 0 73232 0 -1 103360
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3228
timestamp 1644511149
transform 1 0 78384 0 -1 103360
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3229
timestamp 1644511149
transform 1 0 3680 0 1 103360
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3230
timestamp 1644511149
transform 1 0 8832 0 1 103360
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3231
timestamp 1644511149
transform 1 0 13984 0 1 103360
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3232
timestamp 1644511149
transform 1 0 19136 0 1 103360
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3233
timestamp 1644511149
transform 1 0 24288 0 1 103360
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3234
timestamp 1644511149
transform 1 0 29440 0 1 103360
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3235
timestamp 1644511149
transform 1 0 34592 0 1 103360
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3236
timestamp 1644511149
transform 1 0 39744 0 1 103360
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3237
timestamp 1644511149
transform 1 0 44896 0 1 103360
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3238
timestamp 1644511149
transform 1 0 50048 0 1 103360
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3239
timestamp 1644511149
transform 1 0 55200 0 1 103360
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3240
timestamp 1644511149
transform 1 0 60352 0 1 103360
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3241
timestamp 1644511149
transform 1 0 65504 0 1 103360
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3242
timestamp 1644511149
transform 1 0 70656 0 1 103360
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3243
timestamp 1644511149
transform 1 0 75808 0 1 103360
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3244
timestamp 1644511149
transform 1 0 6256 0 -1 104448
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3245
timestamp 1644511149
transform 1 0 11408 0 -1 104448
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3246
timestamp 1644511149
transform 1 0 16560 0 -1 104448
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3247
timestamp 1644511149
transform 1 0 21712 0 -1 104448
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3248
timestamp 1644511149
transform 1 0 26864 0 -1 104448
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3249
timestamp 1644511149
transform 1 0 32016 0 -1 104448
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3250
timestamp 1644511149
transform 1 0 37168 0 -1 104448
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3251
timestamp 1644511149
transform 1 0 42320 0 -1 104448
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3252
timestamp 1644511149
transform 1 0 47472 0 -1 104448
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3253
timestamp 1644511149
transform 1 0 52624 0 -1 104448
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3254
timestamp 1644511149
transform 1 0 57776 0 -1 104448
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3255
timestamp 1644511149
transform 1 0 62928 0 -1 104448
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3256
timestamp 1644511149
transform 1 0 68080 0 -1 104448
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3257
timestamp 1644511149
transform 1 0 73232 0 -1 104448
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3258
timestamp 1644511149
transform 1 0 78384 0 -1 104448
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3259
timestamp 1644511149
transform 1 0 3680 0 1 104448
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3260
timestamp 1644511149
transform 1 0 8832 0 1 104448
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3261
timestamp 1644511149
transform 1 0 13984 0 1 104448
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3262
timestamp 1644511149
transform 1 0 19136 0 1 104448
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3263
timestamp 1644511149
transform 1 0 24288 0 1 104448
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3264
timestamp 1644511149
transform 1 0 29440 0 1 104448
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3265
timestamp 1644511149
transform 1 0 34592 0 1 104448
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3266
timestamp 1644511149
transform 1 0 39744 0 1 104448
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3267
timestamp 1644511149
transform 1 0 44896 0 1 104448
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3268
timestamp 1644511149
transform 1 0 50048 0 1 104448
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3269
timestamp 1644511149
transform 1 0 55200 0 1 104448
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3270
timestamp 1644511149
transform 1 0 60352 0 1 104448
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3271
timestamp 1644511149
transform 1 0 65504 0 1 104448
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3272
timestamp 1644511149
transform 1 0 70656 0 1 104448
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3273
timestamp 1644511149
transform 1 0 75808 0 1 104448
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3274
timestamp 1644511149
transform 1 0 6256 0 -1 105536
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3275
timestamp 1644511149
transform 1 0 11408 0 -1 105536
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3276
timestamp 1644511149
transform 1 0 16560 0 -1 105536
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3277
timestamp 1644511149
transform 1 0 21712 0 -1 105536
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3278
timestamp 1644511149
transform 1 0 26864 0 -1 105536
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3279
timestamp 1644511149
transform 1 0 32016 0 -1 105536
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3280
timestamp 1644511149
transform 1 0 37168 0 -1 105536
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3281
timestamp 1644511149
transform 1 0 42320 0 -1 105536
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3282
timestamp 1644511149
transform 1 0 47472 0 -1 105536
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3283
timestamp 1644511149
transform 1 0 52624 0 -1 105536
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3284
timestamp 1644511149
transform 1 0 57776 0 -1 105536
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3285
timestamp 1644511149
transform 1 0 62928 0 -1 105536
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3286
timestamp 1644511149
transform 1 0 68080 0 -1 105536
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3287
timestamp 1644511149
transform 1 0 73232 0 -1 105536
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3288
timestamp 1644511149
transform 1 0 78384 0 -1 105536
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3289
timestamp 1644511149
transform 1 0 3680 0 1 105536
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3290
timestamp 1644511149
transform 1 0 8832 0 1 105536
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3291
timestamp 1644511149
transform 1 0 13984 0 1 105536
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3292
timestamp 1644511149
transform 1 0 19136 0 1 105536
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3293
timestamp 1644511149
transform 1 0 24288 0 1 105536
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3294
timestamp 1644511149
transform 1 0 29440 0 1 105536
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3295
timestamp 1644511149
transform 1 0 34592 0 1 105536
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3296
timestamp 1644511149
transform 1 0 39744 0 1 105536
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3297
timestamp 1644511149
transform 1 0 44896 0 1 105536
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3298
timestamp 1644511149
transform 1 0 50048 0 1 105536
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3299
timestamp 1644511149
transform 1 0 55200 0 1 105536
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3300
timestamp 1644511149
transform 1 0 60352 0 1 105536
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3301
timestamp 1644511149
transform 1 0 65504 0 1 105536
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3302
timestamp 1644511149
transform 1 0 70656 0 1 105536
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3303
timestamp 1644511149
transform 1 0 75808 0 1 105536
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3304
timestamp 1644511149
transform 1 0 6256 0 -1 106624
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3305
timestamp 1644511149
transform 1 0 11408 0 -1 106624
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3306
timestamp 1644511149
transform 1 0 16560 0 -1 106624
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3307
timestamp 1644511149
transform 1 0 21712 0 -1 106624
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3308
timestamp 1644511149
transform 1 0 26864 0 -1 106624
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3309
timestamp 1644511149
transform 1 0 32016 0 -1 106624
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3310
timestamp 1644511149
transform 1 0 37168 0 -1 106624
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3311
timestamp 1644511149
transform 1 0 42320 0 -1 106624
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3312
timestamp 1644511149
transform 1 0 47472 0 -1 106624
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3313
timestamp 1644511149
transform 1 0 52624 0 -1 106624
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3314
timestamp 1644511149
transform 1 0 57776 0 -1 106624
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3315
timestamp 1644511149
transform 1 0 62928 0 -1 106624
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3316
timestamp 1644511149
transform 1 0 68080 0 -1 106624
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3317
timestamp 1644511149
transform 1 0 73232 0 -1 106624
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3318
timestamp 1644511149
transform 1 0 78384 0 -1 106624
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3319
timestamp 1644511149
transform 1 0 3680 0 1 106624
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3320
timestamp 1644511149
transform 1 0 8832 0 1 106624
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3321
timestamp 1644511149
transform 1 0 13984 0 1 106624
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3322
timestamp 1644511149
transform 1 0 19136 0 1 106624
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3323
timestamp 1644511149
transform 1 0 24288 0 1 106624
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3324
timestamp 1644511149
transform 1 0 29440 0 1 106624
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3325
timestamp 1644511149
transform 1 0 34592 0 1 106624
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3326
timestamp 1644511149
transform 1 0 39744 0 1 106624
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3327
timestamp 1644511149
transform 1 0 44896 0 1 106624
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3328
timestamp 1644511149
transform 1 0 50048 0 1 106624
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3329
timestamp 1644511149
transform 1 0 55200 0 1 106624
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3330
timestamp 1644511149
transform 1 0 60352 0 1 106624
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3331
timestamp 1644511149
transform 1 0 65504 0 1 106624
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3332
timestamp 1644511149
transform 1 0 70656 0 1 106624
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3333
timestamp 1644511149
transform 1 0 75808 0 1 106624
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3334
timestamp 1644511149
transform 1 0 6256 0 -1 107712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3335
timestamp 1644511149
transform 1 0 11408 0 -1 107712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3336
timestamp 1644511149
transform 1 0 16560 0 -1 107712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3337
timestamp 1644511149
transform 1 0 21712 0 -1 107712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3338
timestamp 1644511149
transform 1 0 26864 0 -1 107712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3339
timestamp 1644511149
transform 1 0 32016 0 -1 107712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3340
timestamp 1644511149
transform 1 0 37168 0 -1 107712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3341
timestamp 1644511149
transform 1 0 42320 0 -1 107712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3342
timestamp 1644511149
transform 1 0 47472 0 -1 107712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3343
timestamp 1644511149
transform 1 0 52624 0 -1 107712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3344
timestamp 1644511149
transform 1 0 57776 0 -1 107712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3345
timestamp 1644511149
transform 1 0 62928 0 -1 107712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3346
timestamp 1644511149
transform 1 0 68080 0 -1 107712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3347
timestamp 1644511149
transform 1 0 73232 0 -1 107712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3348
timestamp 1644511149
transform 1 0 78384 0 -1 107712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3349
timestamp 1644511149
transform 1 0 3680 0 1 107712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3350
timestamp 1644511149
transform 1 0 8832 0 1 107712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3351
timestamp 1644511149
transform 1 0 13984 0 1 107712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3352
timestamp 1644511149
transform 1 0 19136 0 1 107712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3353
timestamp 1644511149
transform 1 0 24288 0 1 107712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3354
timestamp 1644511149
transform 1 0 29440 0 1 107712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3355
timestamp 1644511149
transform 1 0 34592 0 1 107712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3356
timestamp 1644511149
transform 1 0 39744 0 1 107712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3357
timestamp 1644511149
transform 1 0 44896 0 1 107712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3358
timestamp 1644511149
transform 1 0 50048 0 1 107712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3359
timestamp 1644511149
transform 1 0 55200 0 1 107712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3360
timestamp 1644511149
transform 1 0 60352 0 1 107712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3361
timestamp 1644511149
transform 1 0 65504 0 1 107712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3362
timestamp 1644511149
transform 1 0 70656 0 1 107712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3363
timestamp 1644511149
transform 1 0 75808 0 1 107712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3364
timestamp 1644511149
transform 1 0 6256 0 -1 108800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3365
timestamp 1644511149
transform 1 0 11408 0 -1 108800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3366
timestamp 1644511149
transform 1 0 16560 0 -1 108800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3367
timestamp 1644511149
transform 1 0 21712 0 -1 108800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3368
timestamp 1644511149
transform 1 0 26864 0 -1 108800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3369
timestamp 1644511149
transform 1 0 32016 0 -1 108800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3370
timestamp 1644511149
transform 1 0 37168 0 -1 108800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3371
timestamp 1644511149
transform 1 0 42320 0 -1 108800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3372
timestamp 1644511149
transform 1 0 47472 0 -1 108800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3373
timestamp 1644511149
transform 1 0 52624 0 -1 108800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3374
timestamp 1644511149
transform 1 0 57776 0 -1 108800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3375
timestamp 1644511149
transform 1 0 62928 0 -1 108800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3376
timestamp 1644511149
transform 1 0 68080 0 -1 108800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3377
timestamp 1644511149
transform 1 0 73232 0 -1 108800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3378
timestamp 1644511149
transform 1 0 78384 0 -1 108800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3379
timestamp 1644511149
transform 1 0 3680 0 1 108800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3380
timestamp 1644511149
transform 1 0 8832 0 1 108800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3381
timestamp 1644511149
transform 1 0 13984 0 1 108800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3382
timestamp 1644511149
transform 1 0 19136 0 1 108800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3383
timestamp 1644511149
transform 1 0 24288 0 1 108800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3384
timestamp 1644511149
transform 1 0 29440 0 1 108800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3385
timestamp 1644511149
transform 1 0 34592 0 1 108800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3386
timestamp 1644511149
transform 1 0 39744 0 1 108800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3387
timestamp 1644511149
transform 1 0 44896 0 1 108800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3388
timestamp 1644511149
transform 1 0 50048 0 1 108800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3389
timestamp 1644511149
transform 1 0 55200 0 1 108800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3390
timestamp 1644511149
transform 1 0 60352 0 1 108800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3391
timestamp 1644511149
transform 1 0 65504 0 1 108800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3392
timestamp 1644511149
transform 1 0 70656 0 1 108800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3393
timestamp 1644511149
transform 1 0 75808 0 1 108800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3394
timestamp 1644511149
transform 1 0 6256 0 -1 109888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3395
timestamp 1644511149
transform 1 0 11408 0 -1 109888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3396
timestamp 1644511149
transform 1 0 16560 0 -1 109888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3397
timestamp 1644511149
transform 1 0 21712 0 -1 109888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3398
timestamp 1644511149
transform 1 0 26864 0 -1 109888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3399
timestamp 1644511149
transform 1 0 32016 0 -1 109888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3400
timestamp 1644511149
transform 1 0 37168 0 -1 109888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3401
timestamp 1644511149
transform 1 0 42320 0 -1 109888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3402
timestamp 1644511149
transform 1 0 47472 0 -1 109888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3403
timestamp 1644511149
transform 1 0 52624 0 -1 109888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3404
timestamp 1644511149
transform 1 0 57776 0 -1 109888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3405
timestamp 1644511149
transform 1 0 62928 0 -1 109888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3406
timestamp 1644511149
transform 1 0 68080 0 -1 109888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3407
timestamp 1644511149
transform 1 0 73232 0 -1 109888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3408
timestamp 1644511149
transform 1 0 78384 0 -1 109888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3409
timestamp 1644511149
transform 1 0 3680 0 1 109888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3410
timestamp 1644511149
transform 1 0 8832 0 1 109888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3411
timestamp 1644511149
transform 1 0 13984 0 1 109888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3412
timestamp 1644511149
transform 1 0 19136 0 1 109888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3413
timestamp 1644511149
transform 1 0 24288 0 1 109888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3414
timestamp 1644511149
transform 1 0 29440 0 1 109888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3415
timestamp 1644511149
transform 1 0 34592 0 1 109888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3416
timestamp 1644511149
transform 1 0 39744 0 1 109888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3417
timestamp 1644511149
transform 1 0 44896 0 1 109888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3418
timestamp 1644511149
transform 1 0 50048 0 1 109888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3419
timestamp 1644511149
transform 1 0 55200 0 1 109888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3420
timestamp 1644511149
transform 1 0 60352 0 1 109888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3421
timestamp 1644511149
transform 1 0 65504 0 1 109888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3422
timestamp 1644511149
transform 1 0 70656 0 1 109888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3423
timestamp 1644511149
transform 1 0 75808 0 1 109888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3424
timestamp 1644511149
transform 1 0 6256 0 -1 110976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3425
timestamp 1644511149
transform 1 0 11408 0 -1 110976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3426
timestamp 1644511149
transform 1 0 16560 0 -1 110976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3427
timestamp 1644511149
transform 1 0 21712 0 -1 110976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3428
timestamp 1644511149
transform 1 0 26864 0 -1 110976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3429
timestamp 1644511149
transform 1 0 32016 0 -1 110976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3430
timestamp 1644511149
transform 1 0 37168 0 -1 110976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3431
timestamp 1644511149
transform 1 0 42320 0 -1 110976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3432
timestamp 1644511149
transform 1 0 47472 0 -1 110976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3433
timestamp 1644511149
transform 1 0 52624 0 -1 110976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3434
timestamp 1644511149
transform 1 0 57776 0 -1 110976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3435
timestamp 1644511149
transform 1 0 62928 0 -1 110976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3436
timestamp 1644511149
transform 1 0 68080 0 -1 110976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3437
timestamp 1644511149
transform 1 0 73232 0 -1 110976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3438
timestamp 1644511149
transform 1 0 78384 0 -1 110976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3439
timestamp 1644511149
transform 1 0 3680 0 1 110976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3440
timestamp 1644511149
transform 1 0 8832 0 1 110976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3441
timestamp 1644511149
transform 1 0 13984 0 1 110976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3442
timestamp 1644511149
transform 1 0 19136 0 1 110976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3443
timestamp 1644511149
transform 1 0 24288 0 1 110976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3444
timestamp 1644511149
transform 1 0 29440 0 1 110976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3445
timestamp 1644511149
transform 1 0 34592 0 1 110976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3446
timestamp 1644511149
transform 1 0 39744 0 1 110976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3447
timestamp 1644511149
transform 1 0 44896 0 1 110976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3448
timestamp 1644511149
transform 1 0 50048 0 1 110976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3449
timestamp 1644511149
transform 1 0 55200 0 1 110976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3450
timestamp 1644511149
transform 1 0 60352 0 1 110976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3451
timestamp 1644511149
transform 1 0 65504 0 1 110976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3452
timestamp 1644511149
transform 1 0 70656 0 1 110976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3453
timestamp 1644511149
transform 1 0 75808 0 1 110976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3454
timestamp 1644511149
transform 1 0 6256 0 -1 112064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3455
timestamp 1644511149
transform 1 0 11408 0 -1 112064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3456
timestamp 1644511149
transform 1 0 16560 0 -1 112064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3457
timestamp 1644511149
transform 1 0 21712 0 -1 112064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3458
timestamp 1644511149
transform 1 0 26864 0 -1 112064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3459
timestamp 1644511149
transform 1 0 32016 0 -1 112064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3460
timestamp 1644511149
transform 1 0 37168 0 -1 112064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3461
timestamp 1644511149
transform 1 0 42320 0 -1 112064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3462
timestamp 1644511149
transform 1 0 47472 0 -1 112064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3463
timestamp 1644511149
transform 1 0 52624 0 -1 112064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3464
timestamp 1644511149
transform 1 0 57776 0 -1 112064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3465
timestamp 1644511149
transform 1 0 62928 0 -1 112064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3466
timestamp 1644511149
transform 1 0 68080 0 -1 112064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3467
timestamp 1644511149
transform 1 0 73232 0 -1 112064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3468
timestamp 1644511149
transform 1 0 78384 0 -1 112064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3469
timestamp 1644511149
transform 1 0 3680 0 1 112064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3470
timestamp 1644511149
transform 1 0 8832 0 1 112064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3471
timestamp 1644511149
transform 1 0 13984 0 1 112064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3472
timestamp 1644511149
transform 1 0 19136 0 1 112064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3473
timestamp 1644511149
transform 1 0 24288 0 1 112064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3474
timestamp 1644511149
transform 1 0 29440 0 1 112064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3475
timestamp 1644511149
transform 1 0 34592 0 1 112064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3476
timestamp 1644511149
transform 1 0 39744 0 1 112064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3477
timestamp 1644511149
transform 1 0 44896 0 1 112064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3478
timestamp 1644511149
transform 1 0 50048 0 1 112064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3479
timestamp 1644511149
transform 1 0 55200 0 1 112064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3480
timestamp 1644511149
transform 1 0 60352 0 1 112064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3481
timestamp 1644511149
transform 1 0 65504 0 1 112064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3482
timestamp 1644511149
transform 1 0 70656 0 1 112064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3483
timestamp 1644511149
transform 1 0 75808 0 1 112064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3484
timestamp 1644511149
transform 1 0 6256 0 -1 113152
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3485
timestamp 1644511149
transform 1 0 11408 0 -1 113152
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3486
timestamp 1644511149
transform 1 0 16560 0 -1 113152
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3487
timestamp 1644511149
transform 1 0 21712 0 -1 113152
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3488
timestamp 1644511149
transform 1 0 26864 0 -1 113152
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3489
timestamp 1644511149
transform 1 0 32016 0 -1 113152
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3490
timestamp 1644511149
transform 1 0 37168 0 -1 113152
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3491
timestamp 1644511149
transform 1 0 42320 0 -1 113152
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3492
timestamp 1644511149
transform 1 0 47472 0 -1 113152
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3493
timestamp 1644511149
transform 1 0 52624 0 -1 113152
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3494
timestamp 1644511149
transform 1 0 57776 0 -1 113152
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3495
timestamp 1644511149
transform 1 0 62928 0 -1 113152
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3496
timestamp 1644511149
transform 1 0 68080 0 -1 113152
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3497
timestamp 1644511149
transform 1 0 73232 0 -1 113152
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3498
timestamp 1644511149
transform 1 0 78384 0 -1 113152
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3499
timestamp 1644511149
transform 1 0 3680 0 1 113152
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3500
timestamp 1644511149
transform 1 0 8832 0 1 113152
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3501
timestamp 1644511149
transform 1 0 13984 0 1 113152
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3502
timestamp 1644511149
transform 1 0 19136 0 1 113152
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3503
timestamp 1644511149
transform 1 0 24288 0 1 113152
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3504
timestamp 1644511149
transform 1 0 29440 0 1 113152
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3505
timestamp 1644511149
transform 1 0 34592 0 1 113152
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3506
timestamp 1644511149
transform 1 0 39744 0 1 113152
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3507
timestamp 1644511149
transform 1 0 44896 0 1 113152
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3508
timestamp 1644511149
transform 1 0 50048 0 1 113152
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3509
timestamp 1644511149
transform 1 0 55200 0 1 113152
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3510
timestamp 1644511149
transform 1 0 60352 0 1 113152
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3511
timestamp 1644511149
transform 1 0 65504 0 1 113152
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3512
timestamp 1644511149
transform 1 0 70656 0 1 113152
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3513
timestamp 1644511149
transform 1 0 75808 0 1 113152
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3514
timestamp 1644511149
transform 1 0 6256 0 -1 114240
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3515
timestamp 1644511149
transform 1 0 11408 0 -1 114240
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3516
timestamp 1644511149
transform 1 0 16560 0 -1 114240
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3517
timestamp 1644511149
transform 1 0 21712 0 -1 114240
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3518
timestamp 1644511149
transform 1 0 26864 0 -1 114240
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3519
timestamp 1644511149
transform 1 0 32016 0 -1 114240
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3520
timestamp 1644511149
transform 1 0 37168 0 -1 114240
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3521
timestamp 1644511149
transform 1 0 42320 0 -1 114240
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3522
timestamp 1644511149
transform 1 0 47472 0 -1 114240
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3523
timestamp 1644511149
transform 1 0 52624 0 -1 114240
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3524
timestamp 1644511149
transform 1 0 57776 0 -1 114240
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3525
timestamp 1644511149
transform 1 0 62928 0 -1 114240
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3526
timestamp 1644511149
transform 1 0 68080 0 -1 114240
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3527
timestamp 1644511149
transform 1 0 73232 0 -1 114240
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3528
timestamp 1644511149
transform 1 0 78384 0 -1 114240
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3529
timestamp 1644511149
transform 1 0 3680 0 1 114240
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3530
timestamp 1644511149
transform 1 0 8832 0 1 114240
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3531
timestamp 1644511149
transform 1 0 13984 0 1 114240
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3532
timestamp 1644511149
transform 1 0 19136 0 1 114240
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3533
timestamp 1644511149
transform 1 0 24288 0 1 114240
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3534
timestamp 1644511149
transform 1 0 29440 0 1 114240
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3535
timestamp 1644511149
transform 1 0 34592 0 1 114240
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3536
timestamp 1644511149
transform 1 0 39744 0 1 114240
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3537
timestamp 1644511149
transform 1 0 44896 0 1 114240
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3538
timestamp 1644511149
transform 1 0 50048 0 1 114240
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3539
timestamp 1644511149
transform 1 0 55200 0 1 114240
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3540
timestamp 1644511149
transform 1 0 60352 0 1 114240
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3541
timestamp 1644511149
transform 1 0 65504 0 1 114240
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3542
timestamp 1644511149
transform 1 0 70656 0 1 114240
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3543
timestamp 1644511149
transform 1 0 75808 0 1 114240
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3544
timestamp 1644511149
transform 1 0 6256 0 -1 115328
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3545
timestamp 1644511149
transform 1 0 11408 0 -1 115328
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3546
timestamp 1644511149
transform 1 0 16560 0 -1 115328
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3547
timestamp 1644511149
transform 1 0 21712 0 -1 115328
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3548
timestamp 1644511149
transform 1 0 26864 0 -1 115328
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3549
timestamp 1644511149
transform 1 0 32016 0 -1 115328
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3550
timestamp 1644511149
transform 1 0 37168 0 -1 115328
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3551
timestamp 1644511149
transform 1 0 42320 0 -1 115328
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3552
timestamp 1644511149
transform 1 0 47472 0 -1 115328
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3553
timestamp 1644511149
transform 1 0 52624 0 -1 115328
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3554
timestamp 1644511149
transform 1 0 57776 0 -1 115328
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3555
timestamp 1644511149
transform 1 0 62928 0 -1 115328
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3556
timestamp 1644511149
transform 1 0 68080 0 -1 115328
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3557
timestamp 1644511149
transform 1 0 73232 0 -1 115328
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3558
timestamp 1644511149
transform 1 0 78384 0 -1 115328
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3559
timestamp 1644511149
transform 1 0 3680 0 1 115328
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3560
timestamp 1644511149
transform 1 0 8832 0 1 115328
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3561
timestamp 1644511149
transform 1 0 13984 0 1 115328
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3562
timestamp 1644511149
transform 1 0 19136 0 1 115328
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3563
timestamp 1644511149
transform 1 0 24288 0 1 115328
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3564
timestamp 1644511149
transform 1 0 29440 0 1 115328
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3565
timestamp 1644511149
transform 1 0 34592 0 1 115328
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3566
timestamp 1644511149
transform 1 0 39744 0 1 115328
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3567
timestamp 1644511149
transform 1 0 44896 0 1 115328
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3568
timestamp 1644511149
transform 1 0 50048 0 1 115328
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3569
timestamp 1644511149
transform 1 0 55200 0 1 115328
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3570
timestamp 1644511149
transform 1 0 60352 0 1 115328
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3571
timestamp 1644511149
transform 1 0 65504 0 1 115328
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3572
timestamp 1644511149
transform 1 0 70656 0 1 115328
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3573
timestamp 1644511149
transform 1 0 75808 0 1 115328
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3574
timestamp 1644511149
transform 1 0 6256 0 -1 116416
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3575
timestamp 1644511149
transform 1 0 11408 0 -1 116416
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3576
timestamp 1644511149
transform 1 0 16560 0 -1 116416
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3577
timestamp 1644511149
transform 1 0 21712 0 -1 116416
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3578
timestamp 1644511149
transform 1 0 26864 0 -1 116416
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3579
timestamp 1644511149
transform 1 0 32016 0 -1 116416
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3580
timestamp 1644511149
transform 1 0 37168 0 -1 116416
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3581
timestamp 1644511149
transform 1 0 42320 0 -1 116416
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3582
timestamp 1644511149
transform 1 0 47472 0 -1 116416
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3583
timestamp 1644511149
transform 1 0 52624 0 -1 116416
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3584
timestamp 1644511149
transform 1 0 57776 0 -1 116416
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3585
timestamp 1644511149
transform 1 0 62928 0 -1 116416
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3586
timestamp 1644511149
transform 1 0 68080 0 -1 116416
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3587
timestamp 1644511149
transform 1 0 73232 0 -1 116416
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3588
timestamp 1644511149
transform 1 0 78384 0 -1 116416
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3589
timestamp 1644511149
transform 1 0 3680 0 1 116416
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3590
timestamp 1644511149
transform 1 0 8832 0 1 116416
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3591
timestamp 1644511149
transform 1 0 13984 0 1 116416
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3592
timestamp 1644511149
transform 1 0 19136 0 1 116416
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3593
timestamp 1644511149
transform 1 0 24288 0 1 116416
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3594
timestamp 1644511149
transform 1 0 29440 0 1 116416
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3595
timestamp 1644511149
transform 1 0 34592 0 1 116416
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3596
timestamp 1644511149
transform 1 0 39744 0 1 116416
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3597
timestamp 1644511149
transform 1 0 44896 0 1 116416
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3598
timestamp 1644511149
transform 1 0 50048 0 1 116416
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3599
timestamp 1644511149
transform 1 0 55200 0 1 116416
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3600
timestamp 1644511149
transform 1 0 60352 0 1 116416
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3601
timestamp 1644511149
transform 1 0 65504 0 1 116416
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3602
timestamp 1644511149
transform 1 0 70656 0 1 116416
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3603
timestamp 1644511149
transform 1 0 75808 0 1 116416
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3604
timestamp 1644511149
transform 1 0 3680 0 -1 117504
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3605
timestamp 1644511149
transform 1 0 6256 0 -1 117504
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3606
timestamp 1644511149
transform 1 0 8832 0 -1 117504
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3607
timestamp 1644511149
transform 1 0 11408 0 -1 117504
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3608
timestamp 1644511149
transform 1 0 13984 0 -1 117504
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3609
timestamp 1644511149
transform 1 0 16560 0 -1 117504
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3610
timestamp 1644511149
transform 1 0 19136 0 -1 117504
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3611
timestamp 1644511149
transform 1 0 21712 0 -1 117504
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3612
timestamp 1644511149
transform 1 0 24288 0 -1 117504
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3613
timestamp 1644511149
transform 1 0 26864 0 -1 117504
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3614
timestamp 1644511149
transform 1 0 29440 0 -1 117504
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3615
timestamp 1644511149
transform 1 0 32016 0 -1 117504
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3616
timestamp 1644511149
transform 1 0 34592 0 -1 117504
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3617
timestamp 1644511149
transform 1 0 37168 0 -1 117504
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3618
timestamp 1644511149
transform 1 0 39744 0 -1 117504
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3619
timestamp 1644511149
transform 1 0 42320 0 -1 117504
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3620
timestamp 1644511149
transform 1 0 44896 0 -1 117504
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3621
timestamp 1644511149
transform 1 0 47472 0 -1 117504
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3622
timestamp 1644511149
transform 1 0 50048 0 -1 117504
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3623
timestamp 1644511149
transform 1 0 52624 0 -1 117504
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3624
timestamp 1644511149
transform 1 0 55200 0 -1 117504
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3625
timestamp 1644511149
transform 1 0 57776 0 -1 117504
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3626
timestamp 1644511149
transform 1 0 60352 0 -1 117504
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3627
timestamp 1644511149
transform 1 0 62928 0 -1 117504
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3628
timestamp 1644511149
transform 1 0 65504 0 -1 117504
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3629
timestamp 1644511149
transform 1 0 68080 0 -1 117504
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3630
timestamp 1644511149
transform 1 0 70656 0 -1 117504
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3631
timestamp 1644511149
transform 1 0 73232 0 -1 117504
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3632
timestamp 1644511149
transform 1 0 75808 0 -1 117504
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_3633
timestamp 1644511149
transform 1 0 78384 0 -1 117504
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _02_ caravel_pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 39468 0 -1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__nand3b_4  _03_ caravel_pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 39928 0 1 64192
box -38 -48 1510 592
use sky130_fd_sc_hd__and3b_1  _04_ caravel_pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 40664 0 -1 65280
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _05_ caravel_pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 40020 0 -1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _06_
timestamp 1644511149
transform 1 0 41308 0 -1 92480
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_4  _07_ caravel_pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 39836 0 1 65280
box -38 -48 2154 592
use sky130_fd_sc_hd__clkbuf_1  _08_
timestamp 1644511149
transform 1 0 2116 0 -1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _09_
timestamp 1644511149
transform 1 0 77832 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _10_ caravel_pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 10488 0 -1 79424
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _11_ caravel_pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 2760 0 1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _12_ caravel_pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 77464 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _13_
timestamp 1644511149
transform 1 0 2668 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _14_ caravel_pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 67804 0 1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _15_
timestamp 1644511149
transform 1 0 1748 0 1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _16_
timestamp 1644511149
transform 1 0 1748 0 1 65280
box -38 -48 406 592
use sky130_fd_sc_hd__buf_6  _17_ caravel_pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 77372 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _18_
timestamp 1644511149
transform 1 0 2576 0 -1 78336
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _19_
timestamp 1644511149
transform 1 0 2760 0 -1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _20_
timestamp 1644511149
transform 1 0 77464 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _21_
timestamp 1644511149
transform 1 0 2668 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _22_
timestamp 1644511149
transform 1 0 76544 0 1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _23_
timestamp 1644511149
transform 1 0 1748 0 1 70720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_6  _24_
timestamp 1644511149
transform 1 0 39836 0 1 59840
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _25_
timestamp 1644511149
transform 1 0 40204 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _26_
timestamp 1644511149
transform -1 0 40388 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _27_
timestamp 1644511149
transform 1 0 40204 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _28_
timestamp 1644511149
transform 1 0 36156 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _29_
timestamp 1644511149
transform 1 0 39836 0 -1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _30_
timestamp 1644511149
transform 1 0 39836 0 -1 89216
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  _31_
timestamp 1644511149
transform 1 0 41032 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _32_
timestamp 1644511149
transform 1 0 66424 0 -1 112064
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _33_
timestamp 1644511149
transform 1 0 62836 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _34_
timestamp 1644511149
transform 1 0 77832 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _35_
timestamp 1644511149
transform 1 0 38824 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _36_
timestamp 1644511149
transform 1 0 77648 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _37_
timestamp 1644511149
transform 1 0 40204 0 1 95744
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _38_
timestamp 1644511149
transform 1 0 41032 0 -1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _39_
timestamp 1644511149
transform 1 0 58420 0 1 100096
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _40_
timestamp 1644511149
transform 1 0 41676 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _41_
timestamp 1644511149
transform 1 0 39836 0 1 108800
box -38 -48 406 592
use sky130_fd_sc_hd__buf_6  _42_
timestamp 1644511149
transform 1 0 39836 0 -1 59840
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _43_
timestamp 1644511149
transform 1 0 14904 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _44_
timestamp 1644511149
transform 1 0 1748 0 1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _45_
timestamp 1644511149
transform 1 0 39836 0 -1 116416
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  _46_
timestamp 1644511149
transform 1 0 39836 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  _47_
timestamp 1644511149
transform 1 0 38916 0 -1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _48_
timestamp 1644511149
transform 1 0 40940 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _49_
timestamp 1644511149
transform 1 0 38088 0 1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _50_
timestamp 1644511149
transform 1 0 74520 0 -1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _51_
timestamp 1644511149
transform 1 0 40572 0 -1 116416
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  _52_
timestamp 1644511149
transform 1 0 39836 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _53_
timestamp 1644511149
transform 1 0 77832 0 1 103360
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _54_
timestamp 1644511149
transform 1 0 19228 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  _55_
timestamp 1644511149
transform 1 0 38916 0 -1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _56_
timestamp 1644511149
transform 1 0 24196 0 -1 114240
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _57_
timestamp 1644511149
transform 1 0 35052 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _58_
timestamp 1644511149
transform 1 0 71576 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _59_
timestamp 1644511149
transform 1 0 40756 0 -1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input1
timestamp 1644511149
transform 1 0 11684 0 -1 117504
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input2
timestamp 1644511149
transform 1 0 1748 0 -1 117504
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input3 caravel_pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 77096 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__buf_4  input4
timestamp 1644511149
transform 1 0 1380 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__buf_8  input5 caravel_pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 63020 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_6  input6
timestamp 1644511149
transform 1 0 7176 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  input7
timestamp 1644511149
transform 1 0 29716 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  input8
timestamp 1644511149
transform 1 0 77464 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input9
timestamp 1644511149
transform 1 0 1380 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  input10
timestamp 1644511149
transform 1 0 70748 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  input11
timestamp 1644511149
transform 1 0 1380 0 1 81600
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1644511149
transform 1 0 77740 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  input13
timestamp 1644511149
transform 1 0 1380 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1644511149
transform 1 0 77740 0 -1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  input15
timestamp 1644511149
transform 1 0 77648 0 1 87040
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  input16
timestamp 1644511149
transform 1 0 77188 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  input17
timestamp 1644511149
transform 1 0 77832 0 1 90304
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 1644511149
transform 1 0 47748 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input19
timestamp 1644511149
transform 1 0 1380 0 1 101184
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input20
timestamp 1644511149
transform 1 0 1748 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input21
timestamp 1644511149
transform 1 0 1380 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input22
timestamp 1644511149
transform 1 0 59064 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_4  input23
timestamp 1644511149
transform 1 0 1748 0 1 116416
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  input24
timestamp 1644511149
transform 1 0 26956 0 -1 117504
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  input25
timestamp 1644511149
transform 1 0 1380 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input26
timestamp 1644511149
transform 1 0 1380 0 -1 97920
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input27
timestamp 1644511149
transform 1 0 14904 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_6  input28
timestamp 1644511149
transform 1 0 3772 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  input29
timestamp 1644511149
transform 1 0 71116 0 -1 117504
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  input30
timestamp 1644511149
transform 1 0 49036 0 -1 117504
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  input31
timestamp 1644511149
transform 1 0 44988 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input32
timestamp 1644511149
transform 1 0 77096 0 -1 117504
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input33
timestamp 1644511149
transform 1 0 77648 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  input34
timestamp 1644511149
transform 1 0 1380 0 1 105536
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input35
timestamp 1644511149
transform 1 0 1748 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input36
timestamp 1644511149
transform 1 0 18124 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input37
timestamp 1644511149
transform 1 0 32936 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input38
timestamp 1644511149
transform 1 0 51612 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input39
timestamp 1644511149
transform 1 0 77464 0 -1 79424
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input40
timestamp 1644511149
transform 1 0 55476 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  input41
timestamp 1644511149
transform 1 0 60444 0 -1 117504
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  input42
timestamp 1644511149
transform 1 0 56120 0 -1 117504
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input43
timestamp 1644511149
transform 1 0 1748 0 -1 109888
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_8  input44 caravel_pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 4600 0 -1 117504
box -38 -48 1050 592
use sky130_fd_sc_hd__buf_2  input45
timestamp 1644511149
transform 1 0 66424 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  input46
timestamp 1644511149
transform 1 0 1380 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  input47
timestamp 1644511149
transform 1 0 1380 0 -1 90304
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  input48
timestamp 1644511149
transform 1 0 77648 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output49
timestamp 1644511149
transform 1 0 1380 0 -1 66368
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output50
timestamp 1644511149
transform 1 0 77648 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output51
timestamp 1644511149
transform 1 0 34684 0 -1 117504
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output52
timestamp 1644511149
transform 1 0 1380 0 -1 94656
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output53
timestamp 1644511149
transform 1 0 77648 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output54
timestamp 1644511149
transform 1 0 1380 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output55
timestamp 1644511149
transform 1 0 45172 0 -1 117504
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output56
timestamp 1644511149
transform 1 0 1380 0 -1 70720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output57
timestamp 1644511149
transform 1 0 1380 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output58
timestamp 1644511149
transform 1 0 77648 0 -1 99008
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output59
timestamp 1644511149
transform 1 0 1380 0 1 78336
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output60
timestamp 1644511149
transform 1 0 1380 0 1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output61
timestamp 1644511149
transform 1 0 77832 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output62
timestamp 1644511149
transform 1 0 1380 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output63
timestamp 1644511149
transform 1 0 77648 0 -1 71808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output64
timestamp 1644511149
transform 1 0 1380 0 1 85952
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output65
timestamp 1644511149
transform -1 0 1748 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output66
timestamp 1644511149
transform 1 0 67068 0 -1 117504
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output67
timestamp 1644511149
transform 1 0 77832 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output68
timestamp 1644511149
transform 1 0 77832 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output69
timestamp 1644511149
transform 1 0 77832 0 1 75072
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output70
timestamp 1644511149
transform 1 0 77648 0 -1 110976
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output71
timestamp 1644511149
transform 1 0 1380 0 1 113152
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output72
timestamp 1644511149
transform 1 0 1380 0 -1 63104
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output73
timestamp 1644511149
transform 1 0 52716 0 -1 117504
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output74
timestamp 1644511149
transform 1 0 40664 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output75
timestamp 1644511149
transform 1 0 74796 0 -1 117504
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output76
timestamp 1644511149
transform 1 0 77832 0 1 114240
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output77
timestamp 1644511149
transform 1 0 21988 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output78
timestamp 1644511149
transform 1 0 11500 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output79
timestamp 1644511149
transform 1 0 1380 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output80
timestamp 1644511149
transform 1 0 77832 0 1 116416
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output81
timestamp 1644511149
transform 1 0 63848 0 -1 117504
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output82
timestamp 1644511149
transform 1 0 77648 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output83
timestamp 1644511149
transform 1 0 74152 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output84
timestamp 1644511149
transform 1 0 77832 0 1 63104
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output85
timestamp 1644511149
transform 1 0 77648 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output86
timestamp 1644511149
transform 1 0 15548 0 -1 117504
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output87
timestamp 1644511149
transform 1 0 19412 0 -1 117504
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output88
timestamp 1644511149
transform 1 0 77832 0 1 94656
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output89
timestamp 1644511149
transform -1 0 1748 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output90
timestamp 1644511149
transform 1 0 25852 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output91
timestamp 1644511149
transform 1 0 77648 0 -1 103360
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output92
timestamp 1644511149
transform 1 0 77832 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output93
timestamp 1644511149
transform 1 0 37444 0 -1 117504
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output94
timestamp 1644511149
transform 1 0 1380 0 1 73984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output95
timestamp 1644511149
transform 1 0 7820 0 -1 117504
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output96
timestamp 1644511149
transform 1 0 22632 0 -1 117504
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output97
timestamp 1644511149
transform 1 0 77648 0 -1 106624
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output98
timestamp 1644511149
transform 1 0 77832 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output99
timestamp 1644511149
transform 1 0 30360 0 -1 117504
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output100
timestamp 1644511149
transform 1 0 37260 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output101
timestamp 1644511149
transform 1 0 77832 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output102
timestamp 1644511149
transform 1 0 77648 0 -1 83776
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output103
timestamp 1644511149
transform -1 0 1748 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output104
timestamp 1644511149
transform 1 0 41308 0 -1 117504
box -38 -48 406 592
<< labels >>
rlabel metal2 s 11610 119200 11666 120000 6 rst_n
port 0 nsew signal input
rlabel metal3 s 0 65968 800 66088 6 sram_addr_a[0]
port 1 nsew signal tristate
rlabel metal3 s 79200 4768 80000 4888 6 sram_addr_a[1]
port 2 nsew signal tristate
rlabel metal2 s 34150 119200 34206 120000 6 sram_addr_a[2]
port 3 nsew signal tristate
rlabel metal3 s 0 93848 800 93968 6 sram_addr_a[3]
port 4 nsew signal tristate
rlabel metal3 s 79200 55768 80000 55888 6 sram_addr_a[4]
port 5 nsew signal tristate
rlabel metal3 s 0 7488 800 7608 6 sram_addr_a[5]
port 6 nsew signal tristate
rlabel metal2 s 45098 119200 45154 120000 6 sram_addr_a[6]
port 7 nsew signal tristate
rlabel metal3 s 0 70048 800 70168 6 sram_addr_a[7]
port 8 nsew signal tristate
rlabel metal3 s 0 34688 800 34808 6 sram_addr_b[0]
port 9 nsew signal tristate
rlabel metal3 s 79200 98608 80000 98728 6 sram_addr_b[1]
port 10 nsew signal tristate
rlabel metal3 s 0 78208 800 78328 6 sram_addr_b[2]
port 11 nsew signal tristate
rlabel metal3 s 0 58488 800 58608 6 sram_addr_b[3]
port 12 nsew signal tristate
rlabel metal3 s 79200 40128 80000 40248 6 sram_addr_b[4]
port 13 nsew signal tristate
rlabel metal3 s 0 46928 800 47048 6 sram_addr_b[5]
port 14 nsew signal tristate
rlabel metal3 s 79200 71408 80000 71528 6 sram_addr_b[6]
port 15 nsew signal tristate
rlabel metal3 s 0 85688 800 85808 6 sram_addr_b[7]
port 16 nsew signal tristate
rlabel metal3 s 0 54408 800 54528 6 sram_csb_a
port 17 nsew signal tristate
rlabel metal2 s 66994 119200 67050 120000 6 sram_csb_b
port 18 nsew signal tristate
rlabel metal3 s 79200 8848 80000 8968 6 sram_din_b[0]
port 19 nsew signal tristate
rlabel metal3 s 79200 36048 80000 36168 6 sram_din_b[10]
port 20 nsew signal tristate
rlabel metal3 s 79200 74808 80000 74928 6 sram_din_b[11]
port 21 nsew signal tristate
rlabel metal3 s 79200 110168 80000 110288 6 sram_din_b[12]
port 22 nsew signal tristate
rlabel metal3 s 0 112888 800 113008 6 sram_din_b[13]
port 23 nsew signal tristate
rlabel metal3 s 0 62568 800 62688 6 sram_din_b[14]
port 24 nsew signal tristate
rlabel metal2 s 52182 119200 52238 120000 6 sram_din_b[15]
port 25 nsew signal tristate
rlabel metal2 s 40590 0 40646 800 6 sram_din_b[16]
port 26 nsew signal tristate
rlabel metal2 s 74722 119200 74778 120000 6 sram_din_b[17]
port 27 nsew signal tristate
rlabel metal3 s 79200 114248 80000 114368 6 sram_din_b[18]
port 28 nsew signal tristate
rlabel metal2 s 21914 0 21970 800 6 sram_din_b[19]
port 29 nsew signal tristate
rlabel metal2 s 10966 0 11022 800 6 sram_din_b[1]
port 30 nsew signal tristate
rlabel metal3 s 0 19048 800 19168 6 sram_din_b[20]
port 31 nsew signal tristate
rlabel metal3 s 79200 118328 80000 118448 6 sram_din_b[21]
port 32 nsew signal tristate
rlabel metal2 s 63774 119200 63830 120000 6 sram_din_b[22]
port 33 nsew signal tristate
rlabel metal3 s 79200 24488 80000 24608 6 sram_din_b[23]
port 34 nsew signal tristate
rlabel metal2 s 74078 0 74134 800 6 sram_din_b[24]
port 35 nsew signal tristate
rlabel metal3 s 79200 63248 80000 63368 6 sram_din_b[25]
port 36 nsew signal tristate
rlabel metal3 s 79200 51688 80000 51808 6 sram_din_b[26]
port 37 nsew signal tristate
rlabel metal2 s 15474 119200 15530 120000 6 sram_din_b[27]
port 38 nsew signal tristate
rlabel metal2 s 19338 119200 19394 120000 6 sram_din_b[28]
port 39 nsew signal tristate
rlabel metal3 s 79200 94528 80000 94648 6 sram_din_b[29]
port 40 nsew signal tristate
rlabel metal3 s 0 15648 800 15768 6 sram_din_b[2]
port 41 nsew signal tristate
rlabel metal2 s 25778 0 25834 800 6 sram_din_b[30]
port 42 nsew signal tristate
rlabel metal3 s 79200 102688 80000 102808 6 sram_din_b[31]
port 43 nsew signal tristate
rlabel metal3 s 79200 20408 80000 20528 6 sram_din_b[3]
port 44 nsew signal tristate
rlabel metal2 s 37370 119200 37426 120000 6 sram_din_b[4]
port 45 nsew signal tristate
rlabel metal3 s 0 74128 800 74248 6 sram_din_b[5]
port 46 nsew signal tristate
rlabel metal2 s 7746 119200 7802 120000 6 sram_din_b[6]
port 47 nsew signal tristate
rlabel metal2 s 22558 119200 22614 120000 6 sram_din_b[7]
port 48 nsew signal tristate
rlabel metal3 s 79200 106088 80000 106208 6 sram_din_b[8]
port 49 nsew signal tristate
rlabel metal3 s 79200 16328 80000 16448 6 sram_din_b[9]
port 50 nsew signal tristate
rlabel metal2 s 30286 119200 30342 120000 6 sram_mask_b[0]
port 51 nsew signal tristate
rlabel metal2 s 36726 0 36782 800 6 sram_mask_b[1]
port 52 nsew signal tristate
rlabel metal3 s 79200 43528 80000 43648 6 sram_mask_b[2]
port 53 nsew signal tristate
rlabel metal3 s 79200 82968 80000 83088 6 sram_mask_b[3]
port 54 nsew signal tristate
rlabel metal3 s 0 50328 800 50448 6 sram_web_b
port 55 nsew signal tristate
rlabel metal5 s 1104 5298 78844 5618 6 vccd1
port 56 nsew power input
rlabel metal5 s 1104 35934 78844 36254 6 vccd1
port 56 nsew power input
rlabel metal5 s 1104 66570 78844 66890 6 vccd1
port 56 nsew power input
rlabel metal5 s 1104 97206 78844 97526 6 vccd1
port 56 nsew power input
rlabel metal4 s 4208 2128 4528 117552 6 vccd1
port 56 nsew power input
rlabel metal4 s 34928 2128 35248 117552 6 vccd1
port 56 nsew power input
rlabel metal4 s 65648 2128 65968 117552 6 vccd1
port 56 nsew power input
rlabel metal5 s 1104 20616 78844 20936 6 vssd1
port 57 nsew ground input
rlabel metal5 s 1104 51252 78844 51572 6 vssd1
port 57 nsew ground input
rlabel metal5 s 1104 81888 78844 82208 6 vssd1
port 57 nsew ground input
rlabel metal5 s 1104 112524 78844 112844 6 vssd1
port 57 nsew ground input
rlabel metal4 s 19568 2128 19888 117552 6 vssd1
port 57 nsew ground input
rlabel metal4 s 50288 2128 50608 117552 6 vssd1
port 57 nsew ground input
rlabel metal2 s 41234 119200 41290 120000 6 wb_ack_o
port 58 nsew signal tristate
rlabel metal2 s 662 119200 718 120000 6 wb_adr_i[0]
port 59 nsew signal input
rlabel metal2 s 77298 0 77354 800 6 wb_adr_i[1]
port 60 nsew signal input
rlabel metal3 s 0 11568 800 11688 6 wb_adr_i[2]
port 61 nsew signal input
rlabel metal2 s 62486 0 62542 800 6 wb_adr_i[3]
port 62 nsew signal input
rlabel metal2 s 7102 0 7158 800 6 wb_adr_i[4]
port 63 nsew signal input
rlabel metal2 s 29642 0 29698 800 6 wb_adr_i[5]
port 64 nsew signal input
rlabel metal3 s 79200 12248 80000 12368 6 wb_adr_i[6]
port 65 nsew signal input
rlabel metal3 s 0 3408 800 3528 6 wb_adr_i[7]
port 66 nsew signal input
rlabel metal3 s 79200 47608 80000 47728 6 wb_clk_i
port 67 nsew signal input
rlabel metal2 s 70214 0 70270 800 6 wb_cyc_i
port 68 nsew signal input
rlabel metal3 s 0 81608 800 81728 6 wb_dat_i[0]
port 69 nsew signal input
rlabel metal3 s 79200 27888 80000 28008 6 wb_dat_i[10]
port 70 nsew signal input
rlabel metal3 s 0 23128 800 23248 6 wb_dat_i[11]
port 71 nsew signal input
rlabel metal3 s 79200 59168 80000 59288 6 wb_dat_i[12]
port 72 nsew signal input
rlabel metal3 s 79200 87048 80000 87168 6 wb_dat_i[13]
port 73 nsew signal input
rlabel metal3 s 79200 688 80000 808 6 wb_dat_i[14]
port 74 nsew signal input
rlabel metal3 s 79200 90448 80000 90568 6 wb_dat_i[15]
port 75 nsew signal input
rlabel metal2 s 47674 0 47730 800 6 wb_dat_i[16]
port 76 nsew signal input
rlabel metal3 s 0 101328 800 101448 6 wb_dat_i[17]
port 77 nsew signal input
rlabel metal3 s 0 42848 800 42968 6 wb_dat_i[18]
port 78 nsew signal input
rlabel metal2 s 18 0 74 800 6 wb_dat_i[19]
port 79 nsew signal input
rlabel metal2 s 59266 0 59322 800 6 wb_dat_i[1]
port 80 nsew signal input
rlabel metal3 s 0 116968 800 117088 6 wb_dat_i[20]
port 81 nsew signal input
rlabel metal2 s 26422 119200 26478 120000 6 wb_dat_i[21]
port 82 nsew signal input
rlabel metal3 s 0 27208 800 27328 6 wb_dat_i[22]
port 83 nsew signal input
rlabel metal3 s 0 97248 800 97368 6 wb_dat_i[23]
port 84 nsew signal input
rlabel metal2 s 14830 0 14886 800 6 wb_dat_i[24]
port 85 nsew signal input
rlabel metal2 s 3238 0 3294 800 6 wb_dat_i[25]
port 86 nsew signal input
rlabel metal2 s 70858 119200 70914 120000 6 wb_dat_i[26]
port 87 nsew signal input
rlabel metal2 s 48962 119200 49018 120000 6 wb_dat_i[27]
port 88 nsew signal input
rlabel metal2 s 44454 0 44510 800 6 wb_dat_i[28]
port 89 nsew signal input
rlabel metal2 s 78586 119200 78642 120000 6 wb_dat_i[29]
port 90 nsew signal input
rlabel metal3 s 79200 31968 80000 32088 6 wb_dat_i[2]
port 91 nsew signal input
rlabel metal3 s 0 105408 800 105528 6 wb_dat_i[30]
port 92 nsew signal input
rlabel metal3 s 0 38768 800 38888 6 wb_dat_i[31]
port 93 nsew signal input
rlabel metal2 s 18050 0 18106 800 6 wb_dat_i[3]
port 94 nsew signal input
rlabel metal2 s 32862 0 32918 800 6 wb_dat_i[4]
port 95 nsew signal input
rlabel metal2 s 51538 0 51594 800 6 wb_dat_i[5]
port 96 nsew signal input
rlabel metal3 s 79200 78888 80000 79008 6 wb_dat_i[6]
port 97 nsew signal input
rlabel metal2 s 55402 0 55458 800 6 wb_dat_i[7]
port 98 nsew signal input
rlabel metal2 s 59910 119200 59966 120000 6 wb_dat_i[8]
port 99 nsew signal input
rlabel metal2 s 56046 119200 56102 120000 6 wb_dat_i[9]
port 100 nsew signal input
rlabel metal3 s 0 109488 800 109608 6 wb_sel_i[0]
port 101 nsew signal input
rlabel metal2 s 4526 119200 4582 120000 6 wb_sel_i[1]
port 102 nsew signal input
rlabel metal2 s 66350 0 66406 800 6 wb_sel_i[2]
port 103 nsew signal input
rlabel metal3 s 0 31288 800 31408 6 wb_sel_i[3]
port 104 nsew signal input
rlabel metal3 s 0 89768 800 89888 6 wb_stb_i
port 105 nsew signal input
rlabel metal3 s 79200 67328 80000 67448 6 wb_we_i
port 106 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 80000 120000
<< end >>
