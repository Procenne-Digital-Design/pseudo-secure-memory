VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO wbuart
  CLASS BLOCK ;
  FOREIGN wbuart ;
  ORIGIN 0.000 0.000 ;
  SIZE 400.000 BY 800.000 ;
  PIN i_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 554.240 400.000 554.840 ;
    END
  END i_clk
  PIN i_cts_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 642.640 400.000 643.240 ;
    END
  END i_cts_n
  PIN i_reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 343.440 4.000 344.040 ;
    END
  END i_reset
  PIN i_uart_rx
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 331.750 796.000 332.030 800.000 ;
    END
  END i_uart_rx
  PIN i_wb_addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 727.640 400.000 728.240 ;
    END
  END i_wb_addr[0]
  PIN i_wb_addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 374.040 4.000 374.640 ;
    END
  END i_wb_addr[1]
  PIN i_wb_cyc
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 700.440 400.000 701.040 ;
    END
  END i_wb_cyc
  PIN i_wb_data[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.030 796.000 87.310 800.000 ;
    END
  END i_wb_data[0]
  PIN i_wb_data[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 496.440 400.000 497.040 ;
    END
  END i_wb_data[10]
  PIN i_wb_data[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.610 0.000 51.890 4.000 ;
    END
  END i_wb_data[11]
  PIN i_wb_data[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 149.640 400.000 150.240 ;
    END
  END i_wb_data[12]
  PIN i_wb_data[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 122.440 400.000 123.040 ;
    END
  END i_wb_data[13]
  PIN i_wb_data[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 295.840 400.000 296.440 ;
    END
  END i_wb_data[14]
  PIN i_wb_data[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 574.640 4.000 575.240 ;
    END
  END i_wb_data[15]
  PIN i_wb_data[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.530 796.000 167.810 800.000 ;
    END
  END i_wb_data[16]
  PIN i_wb_data[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.790 796.000 113.070 800.000 ;
    END
  END i_wb_data[17]
  PIN i_wb_data[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 380.840 400.000 381.440 ;
    END
  END i_wb_data[18]
  PIN i_wb_data[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 459.040 4.000 459.640 ;
    END
  END i_wb_data[19]
  PIN i_wb_data[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 91.840 400.000 92.440 ;
    END
  END i_wb_data[1]
  PIN i_wb_data[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 222.270 796.000 222.550 800.000 ;
    END
  END i_wb_data[20]
  PIN i_wb_data[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 720.840 4.000 721.440 ;
    END
  END i_wb_data[21]
  PIN i_wb_data[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 516.840 4.000 517.440 ;
    END
  END i_wb_data[22]
  PIN i_wb_data[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 584.840 400.000 585.440 ;
    END
  END i_wb_data[23]
  PIN i_wb_data[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 612.040 400.000 612.640 ;
    END
  END i_wb_data[24]
  PIN i_wb_data[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 438.640 400.000 439.240 ;
    END
  END i_wb_data[25]
  PIN i_wb_data[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 207.440 400.000 208.040 ;
    END
  END i_wb_data[26]
  PIN i_wb_data[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 489.640 4.000 490.240 ;
    END
  END i_wb_data[27]
  PIN i_wb_data[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 227.840 4.000 228.440 ;
    END
  END i_wb_data[28]
  PIN i_wb_data[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 386.490 796.000 386.770 800.000 ;
    END
  END i_wb_data[29]
  PIN i_wb_data[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 411.440 400.000 412.040 ;
    END
  END i_wb_data[2]
  PIN i_wb_data[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 112.240 4.000 112.840 ;
    END
  END i_wb_data[30]
  PIN i_wb_data[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 778.640 4.000 779.240 ;
    END
  END i_wb_data[31]
  PIN i_wb_data[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.090 0.000 161.370 4.000 ;
    END
  END i_wb_data[3]
  PIN i_wb_data[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 251.250 796.000 251.530 800.000 ;
    END
  END i_wb_data[4]
  PIN i_wb_data[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 170.040 4.000 170.640 ;
    END
  END i_wb_data[5]
  PIN i_wb_data[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 632.440 4.000 633.040 ;
    END
  END i_wb_data[6]
  PIN i_wb_data[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 141.770 796.000 142.050 800.000 ;
    END
  END i_wb_data[7]
  PIN i_wb_data[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 215.830 0.000 216.110 4.000 ;
    END
  END i_wb_data[8]
  PIN i_wb_data[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 380.050 0.000 380.330 4.000 ;
    END
  END i_wb_data[9]
  PIN i_wb_sel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 669.840 400.000 670.440 ;
    END
  END i_wb_sel[0]
  PIN i_wb_sel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 316.240 4.000 316.840 ;
    END
  END i_wb_sel[1]
  PIN i_wb_sel[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 54.440 4.000 55.040 ;
    END
  END i_wb_sel[2]
  PIN i_wb_sel[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.330 0.000 135.610 4.000 ;
    END
  END i_wb_sel[3]
  PIN i_wb_stb
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 64.640 400.000 65.240 ;
    END
  END i_wb_stb
  PIN i_wb_we
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 353.640 400.000 354.240 ;
    END
  END i_wb_we
  PIN o_rts_n
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 265.240 400.000 265.840 ;
    END
  END o_rts_n
  PIN o_uart_rx_int
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 354.290 0.000 354.570 4.000 ;
    END
  END o_uart_rx_int
  PIN o_uart_rxfifo_int
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 605.240 4.000 605.840 ;
    END
  END o_uart_rxfifo_int
  PIN o_uart_tx
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 180.240 400.000 180.840 ;
    END
  END o_uart_tx
  PIN o_uart_tx_int
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.310 796.000 3.590 800.000 ;
    END
  END o_uart_tx_int
  PIN o_uart_txfifo_int
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 323.040 400.000 323.640 ;
    END
  END o_uart_txfifo_int
  PIN o_wb_ack
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.240 4.000 27.840 ;
    END
  END o_wb_ack
  PIN o_wb_data[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 34.040 400.000 34.640 ;
    END
  END o_wb_data[0]
  PIN o_wb_data[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 401.240 4.000 401.840 ;
    END
  END o_wb_data[10]
  PIN o_wb_data[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 142.840 4.000 143.440 ;
    END
  END o_wb_data[11]
  PIN o_wb_data[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.050 796.000 58.330 800.000 ;
    END
  END o_wb_data[12]
  PIN o_wb_data[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 270.570 0.000 270.850 4.000 ;
    END
  END o_wb_data[13]
  PIN o_wb_data[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END o_wb_data[14]
  PIN o_wb_data[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 258.440 4.000 259.040 ;
    END
  END o_wb_data[15]
  PIN o_wb_data[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.290 796.000 32.570 800.000 ;
    END
  END o_wb_data[16]
  PIN o_wb_data[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.510 796.000 196.790 800.000 ;
    END
  END o_wb_data[17]
  PIN o_wb_data[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 360.730 796.000 361.010 800.000 ;
    END
  END o_wb_data[18]
  PIN o_wb_data[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 431.840 4.000 432.440 ;
    END
  END o_wb_data[19]
  PIN o_wb_data[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.590 0.000 80.870 4.000 ;
    END
  END o_wb_data[1]
  PIN o_wb_data[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.850 0.000 26.130 4.000 ;
    END
  END o_wb_data[20]
  PIN o_wb_data[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 785.440 400.000 786.040 ;
    END
  END o_wb_data[21]
  PIN o_wb_data[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.040 4.000 85.640 ;
    END
  END o_wb_data[22]
  PIN o_wb_data[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 244.810 0.000 245.090 4.000 ;
    END
  END o_wb_data[23]
  PIN o_wb_data[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 758.240 400.000 758.840 ;
    END
  END o_wb_data[24]
  PIN o_wb_data[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 238.040 400.000 238.640 ;
    END
  END o_wb_data[25]
  PIN o_wb_data[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 690.240 4.000 690.840 ;
    END
  END o_wb_data[26]
  PIN o_wb_data[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 285.640 4.000 286.240 ;
    END
  END o_wb_data[27]
  PIN o_wb_data[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.350 0.000 106.630 4.000 ;
    END
  END o_wb_data[28]
  PIN o_wb_data[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.070 0.000 190.350 4.000 ;
    END
  END o_wb_data[29]
  PIN o_wb_data[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 299.550 0.000 299.830 4.000 ;
    END
  END o_wb_data[2]
  PIN o_wb_data[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 527.040 400.000 527.640 ;
    END
  END o_wb_data[30]
  PIN o_wb_data[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 325.310 0.000 325.590 4.000 ;
    END
  END o_wb_data[31]
  PIN o_wb_data[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.990 796.000 306.270 800.000 ;
    END
  END o_wb_data[3]
  PIN o_wb_data[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 277.010 796.000 277.290 800.000 ;
    END
  END o_wb_data[4]
  PIN o_wb_data[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 663.040 4.000 663.640 ;
    END
  END o_wb_data[5]
  PIN o_wb_data[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 748.040 4.000 748.640 ;
    END
  END o_wb_data[6]
  PIN o_wb_data[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 6.840 400.000 7.440 ;
    END
  END o_wb_data[7]
  PIN o_wb_data[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 200.640 4.000 201.240 ;
    END
  END o_wb_data[8]
  PIN o_wb_data[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 547.440 4.000 548.040 ;
    END
  END o_wb_data[9]
  PIN o_wb_stall
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 469.240 400.000 469.840 ;
    END
  END o_wb_stall
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 26.490 394.220 28.090 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.520 179.670 394.220 181.270 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.520 332.850 394.220 334.450 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.520 486.030 394.220 487.630 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.520 639.210 394.220 640.810 ;
    END
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 789.040 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 103.080 394.220 104.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.520 256.260 394.220 257.860 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.520 409.440 394.220 411.040 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.520 562.620 394.220 564.220 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.520 715.800 394.220 717.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 789.040 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 394.220 788.885 ;
      LAYER met1 ;
        RECT 0.070 10.640 394.220 789.040 ;
      LAYER met2 ;
        RECT 0.100 795.720 3.030 796.690 ;
        RECT 3.870 795.720 32.010 796.690 ;
        RECT 32.850 795.720 57.770 796.690 ;
        RECT 58.610 795.720 86.750 796.690 ;
        RECT 87.590 795.720 112.510 796.690 ;
        RECT 113.350 795.720 141.490 796.690 ;
        RECT 142.330 795.720 167.250 796.690 ;
        RECT 168.090 795.720 196.230 796.690 ;
        RECT 197.070 795.720 221.990 796.690 ;
        RECT 222.830 795.720 250.970 796.690 ;
        RECT 251.810 795.720 276.730 796.690 ;
        RECT 277.570 795.720 305.710 796.690 ;
        RECT 306.550 795.720 331.470 796.690 ;
        RECT 332.310 795.720 360.450 796.690 ;
        RECT 361.290 795.720 386.210 796.690 ;
        RECT 387.050 795.720 392.750 796.690 ;
        RECT 0.100 4.280 392.750 795.720 ;
        RECT 0.650 4.000 25.570 4.280 ;
        RECT 26.410 4.000 51.330 4.280 ;
        RECT 52.170 4.000 80.310 4.280 ;
        RECT 81.150 4.000 106.070 4.280 ;
        RECT 106.910 4.000 135.050 4.280 ;
        RECT 135.890 4.000 160.810 4.280 ;
        RECT 161.650 4.000 189.790 4.280 ;
        RECT 190.630 4.000 215.550 4.280 ;
        RECT 216.390 4.000 244.530 4.280 ;
        RECT 245.370 4.000 270.290 4.280 ;
        RECT 271.130 4.000 299.270 4.280 ;
        RECT 300.110 4.000 325.030 4.280 ;
        RECT 325.870 4.000 354.010 4.280 ;
        RECT 354.850 4.000 379.770 4.280 ;
        RECT 380.610 4.000 392.750 4.280 ;
      LAYER met3 ;
        RECT 4.000 786.440 396.000 788.965 ;
        RECT 4.000 785.040 395.600 786.440 ;
        RECT 4.000 779.640 396.000 785.040 ;
        RECT 4.400 778.240 396.000 779.640 ;
        RECT 4.000 759.240 396.000 778.240 ;
        RECT 4.000 757.840 395.600 759.240 ;
        RECT 4.000 749.040 396.000 757.840 ;
        RECT 4.400 747.640 396.000 749.040 ;
        RECT 4.000 728.640 396.000 747.640 ;
        RECT 4.000 727.240 395.600 728.640 ;
        RECT 4.000 721.840 396.000 727.240 ;
        RECT 4.400 720.440 396.000 721.840 ;
        RECT 4.000 701.440 396.000 720.440 ;
        RECT 4.000 700.040 395.600 701.440 ;
        RECT 4.000 691.240 396.000 700.040 ;
        RECT 4.400 689.840 396.000 691.240 ;
        RECT 4.000 670.840 396.000 689.840 ;
        RECT 4.000 669.440 395.600 670.840 ;
        RECT 4.000 664.040 396.000 669.440 ;
        RECT 4.400 662.640 396.000 664.040 ;
        RECT 4.000 643.640 396.000 662.640 ;
        RECT 4.000 642.240 395.600 643.640 ;
        RECT 4.000 633.440 396.000 642.240 ;
        RECT 4.400 632.040 396.000 633.440 ;
        RECT 4.000 613.040 396.000 632.040 ;
        RECT 4.000 611.640 395.600 613.040 ;
        RECT 4.000 606.240 396.000 611.640 ;
        RECT 4.400 604.840 396.000 606.240 ;
        RECT 4.000 585.840 396.000 604.840 ;
        RECT 4.000 584.440 395.600 585.840 ;
        RECT 4.000 575.640 396.000 584.440 ;
        RECT 4.400 574.240 396.000 575.640 ;
        RECT 4.000 555.240 396.000 574.240 ;
        RECT 4.000 553.840 395.600 555.240 ;
        RECT 4.000 548.440 396.000 553.840 ;
        RECT 4.400 547.040 396.000 548.440 ;
        RECT 4.000 528.040 396.000 547.040 ;
        RECT 4.000 526.640 395.600 528.040 ;
        RECT 4.000 517.840 396.000 526.640 ;
        RECT 4.400 516.440 396.000 517.840 ;
        RECT 4.000 497.440 396.000 516.440 ;
        RECT 4.000 496.040 395.600 497.440 ;
        RECT 4.000 490.640 396.000 496.040 ;
        RECT 4.400 489.240 396.000 490.640 ;
        RECT 4.000 470.240 396.000 489.240 ;
        RECT 4.000 468.840 395.600 470.240 ;
        RECT 4.000 460.040 396.000 468.840 ;
        RECT 4.400 458.640 396.000 460.040 ;
        RECT 4.000 439.640 396.000 458.640 ;
        RECT 4.000 438.240 395.600 439.640 ;
        RECT 4.000 432.840 396.000 438.240 ;
        RECT 4.400 431.440 396.000 432.840 ;
        RECT 4.000 412.440 396.000 431.440 ;
        RECT 4.000 411.040 395.600 412.440 ;
        RECT 4.000 402.240 396.000 411.040 ;
        RECT 4.400 400.840 396.000 402.240 ;
        RECT 4.000 381.840 396.000 400.840 ;
        RECT 4.000 380.440 395.600 381.840 ;
        RECT 4.000 375.040 396.000 380.440 ;
        RECT 4.400 373.640 396.000 375.040 ;
        RECT 4.000 354.640 396.000 373.640 ;
        RECT 4.000 353.240 395.600 354.640 ;
        RECT 4.000 344.440 396.000 353.240 ;
        RECT 4.400 343.040 396.000 344.440 ;
        RECT 4.000 324.040 396.000 343.040 ;
        RECT 4.000 322.640 395.600 324.040 ;
        RECT 4.000 317.240 396.000 322.640 ;
        RECT 4.400 315.840 396.000 317.240 ;
        RECT 4.000 296.840 396.000 315.840 ;
        RECT 4.000 295.440 395.600 296.840 ;
        RECT 4.000 286.640 396.000 295.440 ;
        RECT 4.400 285.240 396.000 286.640 ;
        RECT 4.000 266.240 396.000 285.240 ;
        RECT 4.000 264.840 395.600 266.240 ;
        RECT 4.000 259.440 396.000 264.840 ;
        RECT 4.400 258.040 396.000 259.440 ;
        RECT 4.000 239.040 396.000 258.040 ;
        RECT 4.000 237.640 395.600 239.040 ;
        RECT 4.000 228.840 396.000 237.640 ;
        RECT 4.400 227.440 396.000 228.840 ;
        RECT 4.000 208.440 396.000 227.440 ;
        RECT 4.000 207.040 395.600 208.440 ;
        RECT 4.000 201.640 396.000 207.040 ;
        RECT 4.400 200.240 396.000 201.640 ;
        RECT 4.000 181.240 396.000 200.240 ;
        RECT 4.000 179.840 395.600 181.240 ;
        RECT 4.000 171.040 396.000 179.840 ;
        RECT 4.400 169.640 396.000 171.040 ;
        RECT 4.000 150.640 396.000 169.640 ;
        RECT 4.000 149.240 395.600 150.640 ;
        RECT 4.000 143.840 396.000 149.240 ;
        RECT 4.400 142.440 396.000 143.840 ;
        RECT 4.000 123.440 396.000 142.440 ;
        RECT 4.000 122.040 395.600 123.440 ;
        RECT 4.000 113.240 396.000 122.040 ;
        RECT 4.400 111.840 396.000 113.240 ;
        RECT 4.000 92.840 396.000 111.840 ;
        RECT 4.000 91.440 395.600 92.840 ;
        RECT 4.000 86.040 396.000 91.440 ;
        RECT 4.400 84.640 396.000 86.040 ;
        RECT 4.000 65.640 396.000 84.640 ;
        RECT 4.000 64.240 395.600 65.640 ;
        RECT 4.000 55.440 396.000 64.240 ;
        RECT 4.400 54.040 396.000 55.440 ;
        RECT 4.000 35.040 396.000 54.040 ;
        RECT 4.000 33.640 395.600 35.040 ;
        RECT 4.000 28.240 396.000 33.640 ;
        RECT 4.400 26.840 396.000 28.240 ;
        RECT 4.000 7.840 396.000 26.840 ;
        RECT 4.000 6.975 395.600 7.840 ;
      LAYER met4 ;
        RECT 8.575 12.415 20.640 749.185 ;
        RECT 23.040 12.415 97.440 749.185 ;
        RECT 99.840 12.415 174.240 749.185 ;
        RECT 176.640 12.415 248.090 749.185 ;
  END
END wbuart
END LIBRARY

